library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bagman_speech2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bagman_speech2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"C6",X"D4",X"BD",X"9D",X"84",X"94",X"C4",X"C4",X"94",X"84",X"D7",X"8E",X"A4",X"FE",X"C4",
		X"C7",X"BC",X"E5",X"8C",X"AF",X"F6",X"8D",X"8D",X"CF",X"DE",X"A5",X"A6",X"CC",X"95",X"E6",X"EF",
		X"FE",X"94",X"E5",X"94",X"84",X"E5",X"B4",X"97",X"EE",X"E4",X"9F",X"C4",X"85",X"EE",X"F6",X"9E",
		X"ED",X"E7",X"DF",X"EC",X"EC",X"BE",X"85",X"95",X"EE",X"84",X"F7",X"FF",X"DC",X"85",X"F4",X"84",
		X"F5",X"C4",X"B5",X"A7",X"BF",X"B5",X"CE",X"95",X"A5",X"CE",X"C7",X"9E",X"BF",X"87",X"CD",X"BE",
		X"BD",X"B7",X"94",X"ED",X"86",X"DC",X"FE",X"A5",X"8F",X"FC",X"FD",X"84",X"C4",X"C4",X"A5",X"BF",
		X"AE",X"F4",X"B5",X"F7",X"C4",X"D6",X"A7",X"86",X"96",X"C6",X"D4",X"A7",X"86",X"F6",X"85",X"F4",
		X"B4",X"CC",X"A6",X"D4",X"DF",X"D5",X"C5",X"AC",X"EC",X"95",X"B5",X"EE",X"9F",X"B4",X"A4",X"94",
		X"E5",X"EF",X"AF",X"DE",X"AF",X"8E",X"D4",X"F4",X"A6",X"C7",X"B4",X"FC",X"85",X"C5",X"86",X"EC",
		X"F7",X"FD",X"A5",X"AD",X"F4",X"CD",X"D4",X"A6",X"8D",X"9E",X"E7",X"DE",X"ED",X"8F",X"F7",X"86",
		X"F5",X"FE",X"9D",X"A6",X"D5",X"9C",X"F6",X"C6",X"AD",X"BD",X"C7",X"E4",X"8D",X"FD",X"C4",X"95",
		X"85",X"F4",X"BC",X"BE",X"DC",X"AF",X"8E",X"84",X"F4",X"A6",X"C7",X"F6",X"DC",X"A7",X"F5",X"C6",
		X"AD",X"B4",X"E6",X"9E",X"B7",X"FC",X"CD",X"B6",X"EE",X"8D",X"95",X"E4",X"D5",X"EC",X"95",X"DE",
		X"8C",X"F7",X"D6",X"E5",X"A4",X"96",X"D6",X"95",X"D4",X"A7",X"F4",X"84",X"A5",X"A5",X"F7",X"86",
		X"95",X"CE",X"B7",X"B7",X"BF",X"94",X"ED",X"C4",X"9C",X"F4",X"EC",X"9D",X"EE",X"D5",X"A6",X"FC",
		X"C4",X"AE",X"B7",X"AE",X"FF",X"F7",X"FE",X"CE",X"D7",X"A6",X"87",X"BF",X"CF",X"D7",X"E6",X"DF",
		X"F6",X"8E",X"D7",X"F7",X"A7",X"BE",X"C6",X"8E",X"87",X"CE",X"A7",X"FE",X"AE",X"87",X"8F",X"F7",
		X"86",X"9F",X"8F",X"F6",X"F6",X"AE",X"96",X"EF",X"C6",X"FE",X"D6",X"CE",X"9F",X"EE",X"D6",X"A6",
		X"BE",X"C6",X"AF",X"B6",X"AE",X"FF",X"B7",X"FE",X"CF",X"C7",X"B7",X"86",X"BE",X"CE",X"D7",X"E6",
		X"CF",X"D7",X"86",X"FF",X"97",X"AF",X"8E",X"F6",X"FE",X"B6",X"BF",X"86",X"8F",X"F7",X"DE",X"87",
		X"FF",X"C6",X"D7",X"C7",X"B6",X"B7",X"B6",X"D6",X"A7",X"86",X"F6",X"D6",X"C7",X"97",X"E6",X"D6",
		X"A7",X"E6",X"C6",X"A7",X"BE",X"B6",X"C6",X"A7",X"F7",X"C7",X"C6",X"B7",X"8E",X"F7",X"8E",X"96",
		X"A7",X"D6",X"FE",X"87",X"DE",X"FE",X"E6",X"A6",X"D6",X"DF",X"D6",X"9F",X"A6",X"E6",X"D7",X"B7",
		X"AE",X"F7",X"86",X"96",X"87",X"F6",X"B7",X"E7",X"9E",X"E7",X"8E",X"D6",X"F6",X"A7",X"CF",X"B6",
		X"DE",X"AF",X"F6",X"C6",X"A7",X"FE",X"A7",X"FE",X"B7",X"F7",X"C6",X"A7",X"FE",X"87",X"F7",X"87",
		X"96",X"A7",X"D6",X"D6",X"8F",X"D6",X"EE",X"F7",X"A6",X"D7",X"9E",X"86",X"9F",X"AE",X"E7",X"B7",
		X"97",X"86",X"F7",X"9E",X"96",X"DF",X"AF",X"A6",X"EE",X"96",X"E7",X"C6",X"DE",X"FE",X"EF",X"97",
		X"AE",X"F7",X"86",X"C7",X"C6",X"A7",X"F6",X"A7",X"F7",X"F7",X"E7",X"D6",X"D6",X"B6",X"87",X"F7",
		X"87",X"96",X"B7",X"96",X"DF",X"87",X"D6",X"A6",X"C6",X"86",X"F6",X"A7",X"BF",X"A7",X"8E",X"DF",
		X"E7",X"97",X"86",X"DE",X"B7",X"B7",X"DF",X"A7",X"AE",X"F6",X"DE",X"AF",X"9E",X"96",X"E6",X"F7",
		X"9F",X"A6",X"F7",X"86",X"C6",X"E6",X"87",X"D7",X"8F",X"C6",X"BF",X"CE",X"E7",X"F7",X"B6",X"8F",
		X"A7",X"C6",X"CE",X"C7",X"EE",X"F7",X"8E",X"CF",X"EF",X"A7",X"F6",X"86",X"8F",X"97",X"B7",X"87",
		X"D6",X"A7",X"C7",X"86",X"FF",X"D6",X"8E",X"AF",X"C6",X"D7",X"96",X"8E",X"E7",X"86",X"CE",X"E7",
		X"AF",X"87",X"B6",X"FF",X"C6",X"8E",X"FE",X"87",X"8F",X"87",X"EE",X"FF",X"E6",X"C6",X"D7",X"AE",
		X"9F",X"96",X"C7",X"D6",X"C7",X"E6",X"E7",X"86",X"C7",X"B6",X"F7",X"D6",X"B7",X"B6",X"A6",X"E7",
		X"86",X"D7",X"E7",X"9E",X"97",X"E7",X"C6",X"86",X"F7",X"96",X"86",X"9F",X"86",X"E7",X"96",X"CE",
		X"F7",X"AF",X"9F",X"AE",X"EE",X"DF",X"BF",X"9E",X"EF",X"EF",X"AE",X"DE",X"EF",X"CE",X"EF",X"EF",
		X"BE",X"8E",X"BF",X"CF",X"DE",X"FE",X"8F",X"CF",X"8E",X"CF",X"BF",X"EF",X"DE",X"BF",X"BF",X"AF",
		X"EF",X"8E",X"CF",X"FF",X"8E",X"8F",X"CF",X"BE",X"FF",X"BF",X"CE",X"CE",X"CE",X"9E",X"FF",X"8E",
		X"CF",X"FE",X"8F",X"9F",X"EE",X"FE",X"FF",X"AF",X"BE",X"CF",X"CE",X"DE",X"9F",X"AF",X"DE",X"CF",
		X"EE",X"9E",X"AF",X"BE",X"EF",X"DE",X"DF",X"8E",X"EE",X"8F",X"EE",X"BE",X"EF",X"BE",X"DF",X"9E",
		X"EE",X"EF",X"8E",X"EE",X"BF",X"8F",X"BF",X"DF",X"DE",X"BF",X"EE",X"8E",X"BF",X"CE",X"DE",X"AE",
		X"9E",X"CE",X"DE",X"8E",X"FE",X"DE",X"CE",X"8F",X"EF",X"DE",X"AF",X"BF",X"FF",X"9F",X"9F",X"EE",
		X"CF",X"BE",X"CE",X"AF",X"BF",X"EE",X"CE",X"FF",X"CF",X"EE",X"CE",X"AF",X"AE",X"EF",X"8E",X"AF",
		X"EF",X"CE",X"EE",X"AF",X"CF",X"FE",X"8F",X"BE",X"9F",X"CE",X"FE",X"AF",X"CF",X"AF",X"EE",X"9F",
		X"CE",X"BE",X"EE",X"EF",X"FF",X"AF",X"8E",X"CF",X"EF",X"8E",X"8E",X"EF",X"EE",X"8E",X"EE",X"CE",
		X"DF",X"AF",X"DE",X"DE",X"AF",X"EF",X"9E",X"AF",X"8E",X"DE",X"CF",X"FE",X"CF",X"8E",X"EF",X"AF",
		X"8E",X"DF",X"CE",X"EE",X"AF",X"CF",X"8F",X"EE",X"AE",X"9F",X"FE",X"CF",X"BE",X"EF",X"8E",X"DE",
		X"9F",X"DE",X"BE",X"EE",X"EF",X"9F",X"AE",X"DF",X"DE",X"DE",X"AE",X"8E",X"EF",X"DE",X"8E",X"EF",
		X"CE",X"EF",X"8F",X"CF",X"AE",X"9E",X"DF",X"9F",X"BF",X"EE",X"8E",X"DE",X"FE",X"AF",X"DE",X"CF",
		X"AF",X"8E",X"EF",X"DE",X"FE",X"9F",X"EF",X"9F",X"FE",X"8E",X"8F",X"EF",X"EE",X"AF",X"CF",X"AE",
		X"8E",X"8E",X"CF",X"EF",X"8F",X"FE",X"AE",X"FE",X"9F",X"EE",X"CE",X"BF",X"8E",X"FF",X"FE",X"8F",
		X"CF",X"DF",X"DE",X"BF",X"CE",X"8F",X"AF",X"CE",X"BE",X"DE",X"BE",X"BF",X"DE",X"EE",X"AE",X"9E",
		X"8E",X"AE",X"DE",X"BE",X"8E",X"CF",X"AF",X"DE",X"8E",X"DF",X"BF",X"AE",X"DE",X"CE",X"AF",X"8F",
		X"FF",X"CE",X"9F",X"CF",X"EE",X"8E",X"FE",X"AE",X"EF",X"CE",X"FE",X"EE",X"BE",X"8E",X"FE",X"FE",
		X"EE",X"9E",X"8F",X"FF",X"9E",X"8F",X"DE",X"8E",X"FF",X"AF",X"CE",X"8F",X"EE",X"FF",X"AE",X"CE",
		X"CF",X"BE",X"AE",X"DF",X"BE",X"9E",X"FE",X"9E",X"EE",X"8E",X"CE",X"BE",X"AE",X"CF",X"DF",X"EF",
		X"9E",X"BF",X"9F",X"CF",X"9E",X"BF",X"FE",X"FF",X"8E",X"FF",X"FE",X"DE",X"9E",X"EE",X"EF",X"8F",
		X"BF",X"8E",X"BF",X"FE",X"9F",X"9E",X"DF",X"CF",X"AE",X"BE",X"8E",X"8E",X"8E",X"9F",X"BF",X"CE",
		X"CE",X"BF",X"8E",X"AE",X"DF",X"DE",X"9F",X"AF",X"BE",X"8F",X"DE",X"EE",X"DE",X"AE",X"CF",X"DF",
		X"CF",X"FE",X"FF",X"DE",X"8F",X"9F",X"9E",X"8E",X"9F",X"CF",X"AE",X"CF",X"DF",X"FE",X"8E",X"CF",
		X"BF",X"CF",X"EE",X"FF",X"DE",X"DF",X"FF",X"EE",X"DF",X"EE",X"DE",X"EE",X"CE",X"FE",X"EF",X"DE",
		X"CF",X"CE",X"DF",X"CE",X"CF",X"DF",X"FF",X"CE",X"DE",X"FF",X"EE",X"DF",X"DE",X"FF",X"CE",X"CF",
		X"CF",X"FF",X"CE",X"EF",X"CE",X"EF",X"FF",X"DE",X"DE",X"EF",X"FE",X"FF",X"DF",X"DF",X"DE",X"DE",
		X"CF",X"DF",X"EE",X"CE",X"FF",X"FE",X"FF",X"DF",X"EE",X"FF",X"CE",X"FE",X"CE",X"EE",X"DE",X"FF",
		X"DE",X"EE",X"EF",X"FF",X"CE",X"EF",X"FF",X"FF",X"CE",X"DF",X"DE",X"CE",X"DF",X"DF",X"FE",X"CE",
		X"EF",X"EE",X"FF",X"CE",X"EF",X"EE",X"EF",X"FE",X"FF",X"DF",X"CF",X"FE",X"DF",X"FF",X"DF",X"FE",
		X"DE",X"EE",X"FF",X"DE",X"CE",X"DE",X"DE",X"DE",X"DE",X"DE",X"EE",X"CE",X"FF",X"EF",X"DE",X"CF",
		X"EE",X"FF",X"CF",X"CE",X"DF",X"FF",X"EE",X"DE",X"DE",X"EF",X"DF",X"DE",X"CE",X"FE",X"EE",X"DF",
		X"CE",X"CE",X"CE",X"DE",X"CE",X"CE",X"EE",X"CE",X"FF",X"EF",X"FE",X"CE",X"FF",X"DF",X"FF",X"FE",
		X"DF",X"EF",X"FE",X"EF",X"CF",X"EE",X"FF",X"DE",X"DE",X"FE",X"CE",X"EF",X"CE",X"DE",X"CE",X"DE",
		X"CE",X"CE",X"FE",X"CF",X"EF",X"FF",X"DF",X"CE",X"FE",X"FF",X"DE",X"EE",X"DE",X"EF",X"FF",X"EE",
		X"DF",X"EE",X"CE",X"EE",X"DE",X"EE",X"CE",X"DF",X"CE",X"DE",X"CE",X"CE",X"DE",X"CE",X"EE",X"CE",
		X"DF",X"FF",X"FE",X"CE",X"FE",X"CE",X"CF",X"DE",X"DE",X"FF",X"FE",X"CE",X"CE",X"EF",X"DF",X"EF",
		X"DE",X"EE",X"DE",X"DF",X"CE",X"CE",X"DE",X"CE",X"CE",X"DE",X"FE",X"DF",X"DF",X"FF",X"EF",X"DE",
		X"EE",X"DE",X"CE",X"EF",X"CE",X"FE",X"CF",X"EF",X"DE",X"EF",X"FE",X"CF",X"CE",X"DE",X"EE",X"EF",
		X"DE",X"DE",X"DE",X"CE",X"CE",X"DE",X"EF",X"CE",X"DE",X"FE",X"FE",X"CE",X"FE",X"DE",X"CE",X"FF",
		X"CE",X"FE",X"FF",X"CF",X"DE",X"EF",X"EF",X"CE",X"DE",X"DE",X"EE",X"CF",X"DE",X"DE",X"DE",X"CE",
		X"CE",X"DE",X"FE",X"CF",X"CF",X"CF",X"EF",X"DE",X"FE",X"DE",X"CF",X"DE",X"DE",X"EF",X"FE",X"EE",
		X"DE",X"DF",X"FF",X"EE",X"DE",X"CE",X"FE",X"CF",X"CE",X"DE",X"DE",X"DE",X"CE",X"DE",X"EE",X"CF",
		X"DF",X"CE",X"DF",X"DE",X"EE",X"FE",X"CF",X"EE",X"CE",X"FF",X"DE",X"CE",X"DE",X"EF",X"CF",X"DE",
		X"CE",X"CE",X"FE",X"DF",X"CE",X"CE",X"CE",X"CE",X"DE",X"DE",X"DE",X"CE",X"FF",X"FF",X"CF",X"DE",
		X"EE",X"FE",X"FF",X"DE",X"EE",X"DF",X"EE",X"DE",X"CE",X"EF",X"FF",X"DF",X"FE",X"EE",X"EE",X"FF",
		X"CE",X"FE",X"FE",X"EE",X"EE",X"EE",X"FE",X"EF",X"EF",X"EF",X"FF",X"FE",X"EE",X"EE",X"EF",X"EE",
		X"FE",X"FF",X"EE",X"EF",X"EE",X"FF",X"EF",X"FF",X"EE",X"FE",X"FE",X"FF",X"EE",X"FE",X"FE",X"FE",
		X"FE",X"EE",X"EE",X"EF",X"FF",X"EE",X"FE",X"EE",X"FE",X"EE",X"EF",X"FE",X"FE",X"FF",X"EE",X"EE",
		X"FE",X"EF",X"FF",X"FE",X"EE",X"EE",X"EE",X"FF",X"EE",X"EE",X"EE",X"FE",X"FE",X"EE",X"EE",X"FF",
		X"EE",X"FF",X"EF",X"FE",X"EE",X"EE",X"FF",X"FE",X"FE",X"EF",X"FE",X"FE",X"FE",X"EF",X"FF",X"FF",
		X"EE",X"EE",X"FE",X"FF",X"FE",X"FE",X"EE",X"FE",X"FE",X"EE",X"EE",X"EF",X"FF",X"EE",X"EF",X"EE",
		X"FE",X"FF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EE",X"EE",X"FF",X"FE",X"EF",X"EE",X"FE",X"FE",X"EF",
		X"EE",X"EE",X"EE",X"FE",X"EE",X"FE",X"EF",X"EE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"EF",X"EE",
		X"EE",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FF",X"FE",X"FE",
		X"FE",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"94");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
