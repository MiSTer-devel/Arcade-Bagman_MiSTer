library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bagman_sram_8bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(16 downto 0);
	dout : out std_logic_vector(7 downto 0);
	we   : in  std_logic;
	din  : in  std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bagman_sram_8bits is
	type rom is array(0 to  81919) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"00",X"12",X"04",X"03",X"40",X"64",X"06",X"C0",X"40",X"41",X"14",X"9D",X"08",X"24",X"A0",
		X"42",X"06",X"26",X"48",X"18",X"00",X"20",X"40",X"07",X"24",X"0C",X"50",X"01",X"C0",X"04",X"04",
		X"41",X"05",X"01",X"00",X"CC",X"C1",X"60",X"C0",X"29",X"04",X"1C",X"E1",X"08",X"C0",X"01",X"41",
		X"04",X"50",X"02",X"40",X"48",X"C0",X"42",X"2B",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"D9",X"C5",X"D5",X"E5",X"08",X"F5",X"CD",X"47",X"3C",X"AF",X"32",X"00",X"A0",X"F3",X"CD",X"23",
		X"31",X"CD",X"FA",X"38",X"3A",X"42",X"61",X"3C",X"32",X"42",X"61",X"3A",X"74",X"62",X"FE",X"01",
		X"28",X"05",X"3A",X"ED",X"61",X"FE",X"00",X"CC",X"7F",X"0F",X"3A",X"6F",X"62",X"FE",X"01",X"CA",
		X"94",X"03",X"3A",X"10",X"62",X"FE",X"01",X"20",X"22",X"3A",X"54",X"60",X"FE",X"00",X"28",X"1B",
		X"3A",X"F2",X"61",X"FE",X"01",X"28",X"14",X"3A",X"ED",X"61",X"FE",X"01",X"28",X"0D",X"3A",X"82",
		X"65",X"FE",X"E9",X"D2",X"94",X"03",X"FE",X"0F",X"DA",X"94",X"03",X"3A",X"00",X"B8",X"11",X"00",
		X"98",X"21",X"A0",X"65",X"01",X"20",X"00",X"ED",X"B0",X"CD",X"A4",X"34",X"CD",X"3E",X"35",X"3A",
		X"43",X"61",X"3C",X"32",X"43",X"61",X"CD",X"D1",X"10",X"3A",X"6D",X"62",X"3C",X"32",X"6D",X"62",
		X"FD",X"21",X"B8",X"65",X"3A",X"0D",X"60",X"47",X"3A",X"99",X"60",X"B8",X"28",X"05",X"CD",X"CB",
		X"10",X"18",X"0B",X"DD",X"21",X"94",X"65",X"FD",X"21",X"B8",X"65",X"CD",X"01",X"10",X"FD",X"21",
		X"BC",X"65",X"3A",X"0D",X"60",X"47",X"3A",X"9A",X"60",X"B8",X"28",X"05",X"CD",X"CB",X"10",X"18",
		X"0B",X"DD",X"21",X"98",X"65",X"FD",X"21",X"BC",X"65",X"CD",X"01",X"10",X"3A",X"53",X"60",X"FE",
		X"01",X"CA",X"80",X"03",X"CD",X"72",X"04",X"3A",X"51",X"61",X"FE",X"01",X"CA",X"80",X"03",X"CD",
		X"9A",X"5C",X"3A",X"00",X"B8",X"CD",X"F4",X"03",X"CD",X"96",X"2C",X"CD",X"4E",X"34",X"CD",X"D4",
		X"3C",X"3A",X"00",X"B8",X"3A",X"71",X"62",X"32",X"72",X"62",X"3A",X"0C",X"57",X"32",X"71",X"62",
		X"CD",X"FB",X"07",X"3A",X"2C",X"60",X"FE",X"01",X"28",X"06",X"CD",X"84",X"07",X"3A",X"00",X"B8",
		X"CD",X"D5",X"07",X"AF",X"32",X"2C",X"60",X"FD",X"21",X"56",X"61",X"DD",X"21",X"94",X"65",X"11",
		X"48",X"61",X"CD",X"03",X"04",X"FD",X"21",X"57",X"61",X"DD",X"21",X"98",X"65",X"11",X"49",X"61",
		X"CD",X"03",X"04",X"2A",X"38",X"60",X"DD",X"21",X"EB",X"61",X"FD",X"21",X"3A",X"60",X"DD",X"7E",
		X"00",X"DD",X"A6",X"01",X"08",X"11",X"97",X"65",X"3A",X"99",X"60",X"47",X"3A",X"EB",X"61",X"FE",
		X"00",X"C4",X"0E",X"35",X"2A",X"78",X"60",X"DD",X"21",X"EC",X"61",X"FD",X"21",X"7A",X"60",X"11",
		X"9B",X"65",X"3E",X"00",X"08",X"3A",X"9A",X"60",X"47",X"3A",X"EC",X"61",X"FE",X"00",X"C4",X"0E",
		X"35",X"CD",X"B1",X"03",X"3A",X"00",X"B8",X"3A",X"ED",X"61",X"FE",X"00",X"CC",X"83",X"16",X"CD",
		X"9D",X"10",X"3A",X"00",X"B8",X"CD",X"84",X"1D",X"CD",X"84",X"06",X"CD",X"F4",X"31",X"CD",X"D5",
		X"06",X"3A",X"00",X"B8",X"CD",X"B0",X"08",X"CD",X"30",X"08",X"3A",X"00",X"B8",X"CD",X"FF",X"10",
		X"3A",X"ED",X"61",X"FE",X"00",X"CC",X"F4",X"08",X"3A",X"00",X"B8",X"CD",X"3C",X"11",X"3A",X"83",
		X"65",X"F5",X"3D",X"32",X"83",X"65",X"CD",X"5E",X"55",X"F1",X"32",X"83",X"65",X"3A",X"C7",X"61",
		X"FE",X"00",X"CC",X"C7",X"0D",X"3A",X"4E",X"60",X"FE",X"00",X"20",X"22",X"CD",X"5E",X"55",X"CD",
		X"65",X"3D",X"3A",X"14",X"60",X"FE",X"01",X"20",X"07",X"3A",X"12",X"60",X"FE",X"01",X"20",X"0E",
		X"FD",X"21",X"47",X"60",X"DD",X"21",X"80",X"65",X"CD",X"6D",X"0B",X"3A",X"00",X"B8",X"CD",X"10",
		X"10",X"CD",X"4B",X"10",X"3E",X"01",X"32",X"8A",X"62",X"3A",X"0D",X"60",X"32",X"98",X"60",X"21",
		X"14",X"60",X"DD",X"21",X"80",X"65",X"CD",X"27",X"0A",X"3A",X"00",X"B8",X"3A",X"F2",X"61",X"FE",
		X"00",X"20",X"20",X"3A",X"0D",X"60",X"32",X"98",X"60",X"21",X"08",X"60",X"FD",X"21",X"4D",X"60",
		X"DD",X"21",X"80",X"65",X"3A",X"14",X"60",X"4F",X"3A",X"13",X"60",X"06",X"19",X"CD",X"2E",X"0B",
		X"3A",X"00",X"B8",X"3A",X"0D",X"60",X"32",X"98",X"60",X"DD",X"21",X"80",X"65",X"FD",X"21",X"14",
		X"60",X"CD",X"66",X"0A",X"DD",X"21",X"80",X"65",X"21",X"14",X"60",X"CD",X"A0",X"09",X"3A",X"56",
		X"61",X"FE",X"00",X"20",X"35",X"3A",X"11",X"62",X"FE",X"00",X"20",X"11",X"3A",X"3B",X"60",X"FE",
		X"01",X"20",X"07",X"3A",X"12",X"60",X"FE",X"01",X"20",X"03",X"CD",X"6F",X"11",X"FD",X"21",X"57",
		X"60",X"FD",X"22",X"93",X"60",X"2A",X"38",X"60",X"22",X"44",X"60",X"21",X"35",X"60",X"FD",X"21",
		X"27",X"60",X"3A",X"37",X"60",X"FE",X"01",X"C4",X"AD",X"04",X"3A",X"57",X"61",X"FE",X"00",X"20",
		X"3B",X"3A",X"12",X"62",X"FE",X"00",X"20",X"11",X"3A",X"7B",X"60",X"FE",X"01",X"20",X"07",X"3A",
		X"12",X"60",X"FE",X"01",X"20",X"03",X"CD",X"9B",X"11",X"2A",X"78",X"60",X"22",X"44",X"60",X"FD",
		X"21",X"97",X"60",X"FD",X"22",X"93",X"60",X"2A",X"78",X"60",X"22",X"44",X"60",X"21",X"75",X"60",
		X"FD",X"21",X"67",X"60",X"3A",X"77",X"60",X"FE",X"01",X"C4",X"AD",X"04",X"3A",X"9A",X"60",X"32",
		X"98",X"60",X"21",X"7B",X"60",X"DD",X"21",X"98",X"65",X"CD",X"27",X"0A",X"3A",X"00",X"B8",X"3A",
		X"97",X"60",X"3C",X"32",X"97",X"60",X"FD",X"21",X"8F",X"60",X"21",X"77",X"60",X"DD",X"21",X"98",
		X"65",X"3A",X"EC",X"61",X"FE",X"01",X"28",X"12",X"3A",X"9A",X"60",X"32",X"98",X"60",X"3A",X"7B",
		X"60",X"4F",X"3A",X"7A",X"60",X"06",X"26",X"CD",X"2E",X"0B",X"3A",X"99",X"60",X"32",X"98",X"60",
		X"21",X"3B",X"60",X"DD",X"21",X"94",X"65",X"CD",X"27",X"0A",X"3A",X"57",X"60",X"3C",X"32",X"57",
		X"60",X"FD",X"21",X"4F",X"60",X"21",X"37",X"60",X"DD",X"21",X"94",X"65",X"3A",X"EB",X"61",X"FE",
		X"01",X"28",X"12",X"3A",X"99",X"60",X"32",X"98",X"60",X"3A",X"3B",X"60",X"4F",X"3A",X"3A",X"60",
		X"06",X"26",X"CD",X"2E",X"0B",X"3E",X"01",X"32",X"7F",X"62",X"CD",X"C7",X"18",X"3A",X"00",X"B8",
		X"CD",X"F9",X"3D",X"3A",X"F1",X"61",X"FE",X"00",X"CC",X"BC",X"0E",X"CD",X"BE",X"39",X"CD",X"0F",
		X"56",X"CD",X"FD",X"39",X"CD",X"66",X"3C",X"3A",X"00",X"B8",X"3E",X"01",X"32",X"00",X"A0",X"ED",
		X"56",X"F1",X"08",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"FB",
		X"C9",X"3A",X"5E",X"61",X"FE",X"00",X"C8",X"3A",X"0D",X"60",X"FE",X"01",X"20",X"0D",X"3A",X"9F",
		X"65",X"FE",X"80",X"38",X"06",X"3A",X"9E",X"65",X"3D",X"18",X"04",X"3A",X"9E",X"65",X"3C",X"32",
		X"9E",X"65",X"DD",X"21",X"9C",X"65",X"DD",X"35",X"03",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",
		X"32",X"98",X"60",X"CD",X"8C",X"55",X"2A",X"5A",X"61",X"DD",X"21",X"9C",X"65",X"DD",X"34",X"03",
		X"CD",X"0E",X"25",X"C9",X"3A",X"59",X"61",X"FE",X"00",X"C8",X"3A",X"9F",X"65",X"3C",X"3C",X"32",
		X"9F",X"65",X"C9",X"FD",X"7E",X"00",X"FE",X"00",X"C8",X"2A",X"54",X"61",X"3A",X"53",X"61",X"FE",
		X"07",X"20",X"11",X"7E",X"FE",X"FF",X"28",X"14",X"DD",X"77",X"00",X"23",X"22",X"54",X"61",X"AF",
		X"32",X"53",X"61",X"C9",X"3A",X"53",X"61",X"3C",X"32",X"53",X"61",X"C9",X"3E",X"31",X"DD",X"77",
		X"00",X"AF",X"FD",X"77",X"00",X"12",X"C9",X"23",X"22",X"21",X"22",X"23",X"21",X"22",X"23",X"22",
		X"21",X"23",X"21",X"22",X"23",X"21",X"22",X"23",X"21",X"22",X"23",X"22",X"21",X"22",X"23",X"21",
		X"22",X"23",X"22",X"21",X"23",X"21",X"22",X"23",X"21",X"22",X"23",X"21",X"22",X"FF",X"18",X"17",
		X"16",X"15",X"14",X"15",X"14",X"16",X"15",X"16",X"14",X"15",X"14",X"16",X"15",X"14",X"16",X"15",
		X"14",X"FF",X"FD",X"21",X"51",X"61",X"DD",X"21",X"80",X"65",X"2A",X"54",X"61",X"FD",X"7E",X"00",
		X"FE",X"00",X"C8",X"3A",X"53",X"61",X"FE",X"07",X"20",X"11",X"7E",X"FE",X"FF",X"28",X"14",X"DD",
		X"77",X"00",X"23",X"22",X"54",X"61",X"AF",X"32",X"53",X"61",X"C9",X"3A",X"53",X"61",X"3C",X"32",
		X"53",X"61",X"C9",X"3E",X"01",X"32",X"52",X"61",X"C9",X"94",X"65",X"98",X"65",X"FD",X"7E",X"00",
		X"E6",X"10",X"FE",X"10",X"28",X"15",X"FD",X"7E",X"00",X"E6",X"20",X"FE",X"20",X"C0",X"E5",X"2A",
		X"44",X"60",X"7E",X"FE",X"FF",X"E1",X"C0",X"06",X"00",X"18",X"0C",X"E5",X"2A",X"44",X"60",X"2B",
		X"7E",X"FE",X"FF",X"E1",X"C0",X"06",X"80",X"7E",X"FE",X"0B",X"20",X"05",X"3E",X"01",X"77",X"18",
		X"02",X"3C",X"77",X"7E",X"FE",X"01",X"C8",X"FE",X"03",X"C8",X"FE",X"05",X"C8",X"FE",X"08",X"C8",
		X"FE",X"0A",X"CC",X"23",X"05",X"FE",X"02",X"CC",X"23",X"05",X"FE",X"04",X"CC",X"23",X"05",X"FE",
		X"07",X"CC",X"23",X"05",X"FE",X"09",X"CC",X"23",X"05",X"FE",X"06",X"20",X"09",X"3E",X"27",X"DD",
		X"77",X"00",X"CD",X"23",X"05",X"C9",X"FE",X"0B",X"20",X"08",X"3E",X"A7",X"DD",X"77",X"00",X"CD",
		X"23",X"05",X"C9",X"F5",X"C5",X"3A",X"F5",X"61",X"FE",X"00",X"20",X"14",X"3A",X"CF",X"61",X"FE",
		X"00",X"20",X"0D",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"15",X"3F",X"CD",X"18",X"20",
		X"C1",X"F1",X"F5",X"78",X"FE",X"80",X"20",X"14",X"DD",X"7E",X"03",X"3D",X"DD",X"77",X"03",X"AF",
		X"FD",X"2A",X"93",X"60",X"FD",X"77",X"00",X"CD",X"72",X"0F",X"F1",X"C9",X"DD",X"7E",X"03",X"3C",
		X"DD",X"77",X"03",X"AF",X"FD",X"2A",X"93",X"60",X"FD",X"77",X"00",X"CD",X"72",X"0F",X"F1",X"C9",
		X"FD",X"7E",X"00",X"E6",X"80",X"FE",X"80",X"20",X"0F",X"E5",X"2A",X"44",X"60",X"CD",X"FA",X"0C",
		X"E1",X"3A",X"0B",X"60",X"FE",X"02",X"28",X"1A",X"FD",X"7E",X"00",X"E6",X"40",X"FE",X"40",X"C0",
		X"E5",X"2A",X"44",X"60",X"CD",X"69",X"0D",X"E1",X"3A",X"0B",X"60",X"FE",X"02",X"C0",X"06",X"80",
		X"28",X"02",X"06",X"00",X"7E",X"FE",X"0B",X"20",X"05",X"3E",X"01",X"77",X"18",X"02",X"3C",X"77",
		X"7E",X"FE",X"02",X"28",X"2B",X"FE",X"05",X"28",X"27",X"FE",X"09",X"28",X"23",X"FE",X"FF",X"28",
		X"1F",X"FE",X"04",X"CA",X"E0",X"05",X"FE",X"06",X"CC",X"14",X"06",X"FE",X"08",X"CC",X"14",X"06",
		X"FE",X"0A",X"CC",X"14",X"06",X"FE",X"01",X"20",X"19",X"3E",X"31",X"B0",X"DD",X"77",X"00",X"C9",
		X"F5",X"C5",X"47",X"3A",X"64",X"61",X"B8",X"30",X"03",X"C1",X"F1",X"C9",X"C1",X"F1",X"CD",X"14",
		X"06",X"C9",X"FE",X"03",X"20",X"07",X"3E",X"30",X"B0",X"DD",X"77",X"00",X"C9",X"FE",X"07",X"20",
		X"07",X"3E",X"2E",X"B0",X"DD",X"77",X"00",X"C9",X"FE",X"FF",X"20",X"07",X"3E",X"30",X"B0",X"DD",
		X"77",X"00",X"C9",X"C9",X"F5",X"C5",X"3A",X"F5",X"61",X"FE",X"00",X"20",X"14",X"3A",X"CF",X"61",
		X"FE",X"00",X"20",X"0D",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"39",X"3F",X"CD",X"18",
		X"20",X"C1",X"AF",X"FD",X"2A",X"93",X"60",X"FD",X"77",X"00",X"78",X"FE",X"80",X"28",X"19",X"DD",
		X"7E",X"02",X"3C",X"DD",X"77",X"02",X"FE",X"F0",X"20",X"0C",X"3E",X"01",X"DD",X"77",X"02",X"3A",
		X"98",X"60",X"3C",X"32",X"98",X"60",X"F1",X"C9",X"DD",X"7E",X"02",X"3D",X"DD",X"77",X"02",X"FE",
		X"01",X"20",X"0C",X"3E",X"F0",X"DD",X"77",X"02",X"3A",X"98",X"60",X"3D",X"32",X"98",X"60",X"AF",
		X"FD",X"2A",X"93",X"60",X"FD",X"77",X"00",X"F1",X"C9",X"AF",X"32",X"1C",X"60",X"32",X"1D",X"60",
		X"32",X"1E",X"60",X"C9",X"21",X"1C",X"60",X"DD",X"21",X"8A",X"65",X"FD",X"21",X"82",X"65",X"11",
		X"04",X"00",X"7E",X"FE",X"01",X"28",X"0F",X"23",X"DD",X"19",X"7E",X"FE",X"01",X"28",X"07",X"23",
		X"DD",X"19",X"7E",X"FE",X"01",X"C0",X"3E",X"01",X"32",X"30",X"60",X"3A",X"26",X"60",X"E6",X"08",
		X"FE",X"08",X"CC",X"C9",X"06",X"3A",X"26",X"60",X"E6",X"10",X"FE",X"10",X"CC",X"CF",X"06",X"3E",
		X"01",X"32",X"29",X"60",X"3D",X"32",X"2F",X"60",X"C9",X"3E",X"01",X"32",X"2D",X"60",X"C9",X"3E",
		X"01",X"32",X"2E",X"60",X"C9",X"3A",X"30",X"60",X"FE",X"01",X"C0",X"3A",X"2D",X"60",X"FE",X"01",
		X"CC",X"10",X"07",X"3A",X"2E",X"60",X"FE",X"01",X"CC",X"20",X"07",X"3A",X"2F",X"60",X"3C",X"FE",
		X"04",X"28",X"04",X"32",X"2F",X"60",X"C9",X"AF",X"32",X"2D",X"60",X"32",X"2E",X"60",X"32",X"30",
		X"60",X"32",X"29",X"60",X"32",X"25",X"60",X"CD",X"79",X"06",X"3E",X"20",X"32",X"80",X"65",X"C9",
		X"CD",X"30",X"07",X"CD",X"70",X"07",X"FD",X"7E",X"00",X"3D",X"3D",X"3D",X"FD",X"77",X"00",X"C9",
		X"CD",X"30",X"07",X"CD",X"53",X"07",X"FD",X"7E",X"00",X"3C",X"3C",X"3C",X"FD",X"77",X"00",X"C9",
		X"11",X"4F",X"07",X"3A",X"2F",X"60",X"FE",X"04",X"C8",X"83",X"5F",X"7A",X"CE",X"00",X"57",X"1A",
		X"47",X"3A",X"80",X"65",X"E6",X"08",X"B0",X"32",X"80",X"65",X"AF",X"32",X"25",X"60",X"C9",X"1D",
		X"1D",X"1D",X"1D",X"06",X"20",X"C5",X"2A",X"09",X"60",X"CD",X"FA",X"0C",X"3A",X"0B",X"60",X"FE",
		X"02",X"20",X"02",X"C1",X"C9",X"3E",X"01",X"32",X"25",X"60",X"3D",X"32",X"29",X"60",X"C1",X"C9",
		X"06",X"20",X"C5",X"2A",X"09",X"60",X"CD",X"69",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"20",X"E5",
		X"C1",X"10",X"EF",X"C9",X"CD",X"5E",X"55",X"2A",X"09",X"60",X"2B",X"2B",X"2B",X"7E",X"FE",X"DC",
		X"28",X"03",X"FE",X"0B",X"C0",X"3A",X"2A",X"60",X"FE",X"01",X"C8",X"3E",X"01",X"21",X"1E",X"60",
		X"01",X"03",X"00",X"ED",X"B9",X"C8",X"3A",X"26",X"60",X"E6",X"80",X"FE",X"80",X"C0",X"3A",X"54",
		X"60",X"FE",X"00",X"28",X"08",X"3A",X"50",X"60",X"E6",X"80",X"FE",X"80",X"C8",X"3E",X"01",X"32",
		X"28",X"60",X"32",X"2A",X"60",X"3D",X"32",X"2B",X"60",X"3E",X"01",X"32",X"75",X"62",X"21",X"FD",
		X"3E",X"CD",X"18",X"20",X"C9",X"3A",X"2A",X"60",X"FE",X"01",X"C0",X"11",X"F6",X"07",X"3A",X"2B",
		X"60",X"FE",X"05",X"C8",X"83",X"5F",X"7A",X"CE",X"00",X"57",X"1A",X"32",X"80",X"65",X"3A",X"2B",
		X"60",X"3C",X"32",X"2B",X"60",X"C9",X"1C",X"1C",X"1C",X"1C",X"1B",X"3A",X"2A",X"60",X"FE",X"01",
		X"C0",X"3A",X"26",X"60",X"E6",X"80",X"FE",X"80",X"C0",X"3A",X"54",X"60",X"FE",X"00",X"28",X"08",
		X"3A",X"50",X"60",X"E6",X"80",X"FE",X"80",X"C8",X"AF",X"32",X"2A",X"60",X"32",X"28",X"60",X"32",
		X"29",X"60",X"32",X"2B",X"60",X"3E",X"19",X"32",X"80",X"65",X"3E",X"01",X"32",X"2C",X"60",X"C9",
		X"3A",X"2A",X"60",X"FE",X"01",X"C8",X"3A",X"25",X"60",X"FE",X"01",X"C8",X"3A",X"83",X"65",X"3C",
		X"DD",X"21",X"8A",X"65",X"FD",X"21",X"1C",X"60",X"11",X"04",X"00",X"CD",X"5D",X"08",X"DD",X"19",
		X"FD",X"23",X"CD",X"5D",X"08",X"DD",X"19",X"FD",X"23",X"CD",X"5D",X"08",X"C9",X"DD",X"BE",X"01",
		X"20",X"47",X"F5",X"06",X"08",X"3A",X"82",X"65",X"D6",X"05",X"3C",X"F5",X"DD",X"BE",X"00",X"28",
		X"2F",X"F1",X"10",X"F6",X"18",X"2D",X"FD",X"7E",X"00",X"FE",X"00",X"20",X"17",X"E5",X"DD",X"E5",
		X"21",X"00",X"01",X"CD",X"90",X"5C",X"21",X"03",X"3F",X"CD",X"18",X"20",X"3E",X"01",X"32",X"75",
		X"62",X"DD",X"E1",X"E1",X"3E",X"01",X"FD",X"77",X"00",X"3E",X"1A",X"32",X"80",X"65",X"F1",X"C9",
		X"F1",X"18",X"D3",X"AF",X"FD",X"77",X"00",X"F1",X"C9",X"F5",X"AF",X"FD",X"77",X"00",X"F1",X"C9",
		X"DD",X"21",X"19",X"60",X"FD",X"21",X"8B",X"65",X"3E",X"E1",X"08",X"CD",X"DF",X"08",X"DD",X"23",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"3E",X"41",X"08",X"CD",X"DF",X"08",X"DD",X"23",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"3E",X"C9",X"08",X"CD",X"DF",X"08",X"C9",X"3A",
		X"0D",X"60",X"3D",X"DD",X"BE",X"00",X"C2",X"EE",X"08",X"08",X"FD",X"77",X"00",X"C9",X"3E",X"FF",
		X"FD",X"77",X"00",X"C9",X"DD",X"21",X"16",X"60",X"FD",X"21",X"94",X"09",X"21",X"8A",X"65",X"CD",
		X"25",X"09",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"23",X"23",X"23",X"23",
		X"CD",X"25",X"09",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"23",X"23",X"23",
		X"23",X"CD",X"25",X"09",X"C9",X"DD",X"7E",X"00",X"FE",X"00",X"C2",X"61",X"09",X"7E",X"3D",X"77",
		X"F5",X"DD",X"7E",X"06",X"FE",X"00",X"28",X"07",X"3A",X"82",X"65",X"3D",X"32",X"82",X"65",X"F1",
		X"FD",X"BE",X"02",X"CA",X"4C",X"09",X"FE",X"00",X"CA",X"59",X"09",X"C9",X"DD",X"7E",X"03",X"FD",
		X"BE",X"03",X"C0",X"3E",X"01",X"DD",X"77",X"00",X"C9",X"DD",X"7E",X"03",X"3D",X"DD",X"77",X"03",
		X"C9",X"7E",X"3C",X"77",X"F5",X"DD",X"7E",X"06",X"FE",X"00",X"28",X"07",X"3A",X"82",X"65",X"3C",
		X"32",X"82",X"65",X"F1",X"FD",X"BE",X"00",X"CA",X"7F",X"09",X"FE",X"FF",X"28",X"0E",X"C9",X"DD",
		X"7E",X"03",X"FD",X"BE",X"01",X"C0",X"3E",X"00",X"DD",X"77",X"00",X"C9",X"DD",X"7E",X"03",X"3C",
		X"DD",X"77",X"03",X"C9",X"CF",X"01",X"20",X"00",X"80",X"01",X"50",X"00",X"D0",X"02",X"CA",X"01",
		X"3A",X"12",X"60",X"FE",X"00",X"C8",X"3A",X"11",X"60",X"3C",X"32",X"11",X"60",X"FE",X"5F",X"C0",
		X"AF",X"32",X"11",X"60",X"32",X"12",X"60",X"3C",X"32",X"15",X"60",X"3A",X"0D",X"60",X"FE",X"02",
		X"28",X"06",X"FD",X"21",X"E8",X"09",X"18",X"04",X"FD",X"21",X"DF",X"09",X"06",X"09",X"DD",X"7E",
		X"02",X"FD",X"BE",X"00",X"28",X"1B",X"FD",X"23",X"10",X"F4",X"AF",X"77",X"2B",X"77",X"C9",X"94",
		X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",
		X"34",X"3A",X"87",X"65",X"D6",X"00",X"DD",X"BE",X"03",X"28",X"0E",X"D6",X"01",X"DD",X"BE",X"03",
		X"28",X"07",X"C6",X"02",X"DD",X"BE",X"03",X"20",X"D1",X"3A",X"98",X"60",X"FE",X"01",X"28",X"CA",
		X"3A",X"4E",X"60",X"FE",X"00",X"28",X"0A",X"7D",X"FE",X"14",X"20",X"05",X"3E",X"01",X"32",X"25",
		X"60",X"3E",X"01",X"77",X"2B",X"77",X"C9",X"3A",X"98",X"60",X"FE",X"02",X"20",X"06",X"FD",X"21",
		X"42",X"0A",X"18",X"04",X"FD",X"21",X"54",X"0A",X"06",X"12",X"7E",X"F5",X"CD",X"CE",X"09",X"F1",
		X"77",X"C9",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",
		X"9D",X"9E",X"9F",X"A0",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",
		X"33",X"34",X"35",X"36",X"37",X"38",X"3A",X"12",X"60",X"FE",X"00",X"C0",X"21",X"87",X"65",X"3A",
		X"10",X"60",X"FE",X"01",X"20",X"71",X"7E",X"FE",X"12",X"38",X"62",X"3A",X"15",X"60",X"FE",X"01",
		X"CA",X"AE",X"0A",X"3A",X"0D",X"60",X"FE",X"03",X"CA",X"99",X"0A",X"7E",X"FE",X"42",X"CA",X"28",
		X"0B",X"FE",X"6A",X"CA",X"28",X"0B",X"C3",X"AE",X"0A",X"7E",X"FE",X"AA",X"CA",X"28",X"0B",X"FE",
		X"8A",X"CA",X"28",X"0B",X"FE",X"72",X"CA",X"28",X"0B",X"FE",X"2A",X"CA",X"28",X"0B",X"35",X"AF",
		X"32",X"15",X"60",X"FD",X"7E",X"00",X"FE",X"01",X"20",X"07",X"DD",X"7E",X"03",X"3D",X"DD",X"77",
		X"03",X"FD",X"7E",X"27",X"FE",X"01",X"20",X"07",X"DD",X"7E",X"17",X"3D",X"DD",X"77",X"17",X"FD",
		X"7E",X"67",X"FE",X"01",X"C0",X"DD",X"7E",X"1B",X"3D",X"DD",X"77",X"1B",X"C9",X"3E",X"00",X"32",
		X"10",X"60",X"3C",X"32",X"12",X"60",X"C9",X"3A",X"0D",X"60",X"FE",X"03",X"28",X"05",X"7E",X"FE",
		X"89",X"18",X"03",X"7E",X"FE",X"C9",X"30",X"2B",X"34",X"FD",X"7E",X"00",X"FE",X"01",X"20",X"07",
		X"DD",X"7E",X"03",X"3C",X"DD",X"77",X"03",X"FD",X"7E",X"27",X"FE",X"01",X"20",X"07",X"DD",X"7E",
		X"17",X"3C",X"DD",X"77",X"17",X"FD",X"7E",X"67",X"FE",X"01",X"C0",X"DD",X"7E",X"1B",X"3C",X"DD",
		X"77",X"1B",X"C9",X"3E",X"01",X"32",X"10",X"60",X"3E",X"01",X"32",X"12",X"60",X"C9",X"FE",X"01",
		X"28",X"2D",X"7E",X"FE",X"00",X"28",X"28",X"79",X"FE",X"00",X"C0",X"78",X"DD",X"77",X"00",X"DD",
		X"34",X"03",X"FD",X"34",X"00",X"3A",X"F5",X"61",X"FE",X"00",X"C0",X"3E",X"0D",X"47",X"3A",X"98",
		X"60",X"B8",X"C0",X"3E",X"01",X"32",X"F5",X"61",X"21",X"45",X"3F",X"CD",X"18",X"20",X"C9",X"AF",
		X"FD",X"77",X"00",X"C9",X"F1",X"AF",X"32",X"9B",X"60",X"FD",X"77",X"00",X"C9",X"3A",X"25",X"60",
		X"FE",X"01",X"C8",X"3A",X"28",X"60",X"FE",X"01",X"CA",X"65",X"0B",X"3A",X"26",X"60",X"E6",X"10",
		X"FE",X"10",X"20",X"0D",X"2A",X"09",X"60",X"CD",X"FA",X"0C",X"3A",X"0B",X"60",X"FE",X"02",X"28",
		X"1C",X"3A",X"26",X"60",X"E6",X"08",X"FE",X"08",X"C2",X"65",X"0B",X"2A",X"09",X"60",X"CD",X"69",
		X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"C2",X"65",X"0B",X"06",X"80",X"28",X"02",X"06",X"00",X"3A",
		X"06",X"60",X"FE",X"0B",X"20",X"1A",X"3E",X"01",X"32",X"06",X"60",X"C5",X"CD",X"FD",X"0F",X"E5",
		X"DD",X"E5",X"D5",X"21",X"10",X"00",X"CD",X"90",X"5C",X"D1",X"DD",X"E1",X"E1",X"C1",X"18",X"14",
		X"3C",X"F5",X"3A",X"58",X"61",X"FE",X"00",X"28",X"07",X"CD",X"D9",X"0C",X"FE",X"00",X"28",X"39",
		X"F1",X"32",X"06",X"60",X"3A",X"06",X"60",X"21",X"80",X"65",X"FE",X"02",X"CC",X"36",X"0C",X"FE",
		X"05",X"CC",X"36",X"0C",X"FE",X"09",X"CC",X"36",X"0C",X"FE",X"FF",X"C8",X"FE",X"04",X"CC",X"36",
		X"0C",X"FE",X"06",X"CC",X"36",X"0C",X"FE",X"08",X"CC",X"36",X"0C",X"FE",X"0A",X"CC",X"36",X"0C",
		X"FE",X"01",X"20",X"07",X"3E",X"20",X"B0",X"77",X"C9",X"F1",X"C9",X"FE",X"03",X"20",X"05",X"3E",
		X"1F",X"B0",X"77",X"C9",X"FE",X"07",X"20",X"05",X"3E",X"1E",X"B0",X"77",X"C9",X"FE",X"FF",X"20",
		X"04",X"3E",X"80",X"77",X"C9",X"C9",X"F5",X"78",X"FE",X"80",X"28",X"5A",X"2A",X"09",X"60",X"CD",
		X"FA",X"0C",X"3A",X"0B",X"60",X"FE",X"02",X"C2",X"64",X"0B",X"3A",X"82",X"65",X"3C",X"32",X"82",
		X"65",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"1A",X"CD",X"7C",X"0C",X"3A",X"F3",X"61",X"FE",X"00",
		X"20",X"10",X"CD",X"89",X"0C",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"33",X"3F",X"CD",
		X"18",X"20",X"3E",X"01",X"FD",X"77",X"00",X"32",X"9B",X"60",X"F1",X"C9",X"3A",X"CF",X"61",X"FE",
		X"00",X"C8",X"21",X"2D",X"3F",X"CD",X"18",X"20",X"C9",X"3A",X"C7",X"61",X"FE",X"00",X"C9",X"21",
		X"3F",X"3F",X"CD",X"18",X"20",X"C9",X"2A",X"09",X"60",X"CD",X"69",X"0D",X"3A",X"0B",X"60",X"FE",
		X"02",X"C2",X"64",X"0B",X"3A",X"82",X"65",X"3D",X"32",X"82",X"65",X"CD",X"17",X"25",X"3A",X"F3",
		X"61",X"FE",X"00",X"20",X"1A",X"CD",X"7C",X"0C",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"10",X"CD",
		X"89",X"0C",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"33",X"3F",X"CD",X"18",X"20",X"3E",
		X"01",X"FD",X"77",X"00",X"32",X"9B",X"60",X"F1",X"C9",X"C5",X"06",X"02",X"3A",X"7C",X"62",X"FE",
		X"00",X"28",X"02",X"06",X"01",X"3A",X"5F",X"61",X"B8",X"C1",X"38",X"07",X"AF",X"32",X"5F",X"61",
		X"3E",X"00",X"C9",X"3C",X"32",X"5F",X"61",X"3E",X"01",X"C9",X"3A",X"ED",X"61",X"FE",X"01",X"20",
		X"06",X"3E",X"02",X"32",X"0B",X"60",X"C9",X"3A",X"F2",X"61",X"FE",X"01",X"28",X"F3",X"CD",X"85",
		X"25",X"3A",X"0B",X"60",X"FE",X"02",X"C8",X"7D",X"D6",X"21",X"6F",X"7C",X"DE",X"00",X"67",X"7E",
		X"CD",X"A2",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"C0",X"2B",X"7E",X"CD",X"A2",X"0D",X"23",X"23",
		X"CD",X"34",X"0D",X"C9",X"7E",X"E5",X"C5",X"01",X"0D",X"00",X"21",X"45",X"0D",X"ED",X"B1",X"C1",
		X"E1",X"CA",X"52",X"0D",X"C9",X"FB",X"FA",X"BA",X"A4",X"6C",X"66",X"62",X"25",X"22",X"26",X"6D",
		X"78",X"B1",X"DD",X"E5",X"CD",X"40",X"26",X"DD",X"E1",X"78",X"FE",X"05",X"D8",X"3E",X"01",X"32",
		X"0B",X"60",X"C9",X"3E",X"01",X"32",X"0B",X"60",X"C9",X"3A",X"ED",X"61",X"FE",X"01",X"20",X"06",
		X"3E",X"02",X"32",X"0B",X"60",X"C9",X"CD",X"69",X"25",X"3A",X"0B",X"60",X"FE",X"02",X"C8",X"7D",
		X"C6",X"1F",X"6F",X"7C",X"CE",X"00",X"67",X"7E",X"CD",X"A2",X"0D",X"3A",X"0B",X"60",X"FE",X"02",
		X"C0",X"2B",X"7E",X"CD",X"A2",X"0D",X"23",X"23",X"CD",X"34",X"0D",X"C9",X"3E",X"02",X"32",X"0B",
		X"60",X"C9",X"4F",X"11",X"B1",X"0D",X"06",X"16",X"1A",X"B9",X"28",X"F0",X"13",X"10",X"F9",X"18",
		X"B2",X"E0",X"FF",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F0",X"EF",X"EE",X"ED",X"EC",X"EB",X"EA",
		X"F7",X"DF",X"DE",X"DE",X"4B",X"4A",X"49",X"3A",X"9B",X"60",X"FE",X"01",X"C8",X"3A",X"26",X"60",
		X"E6",X"20",X"FE",X"20",X"28",X"13",X"3A",X"26",X"60",X"E6",X"40",X"FE",X"40",X"C0",X"2A",X"09",
		X"60",X"7E",X"FE",X"FF",X"C0",X"06",X"00",X"18",X"0A",X"2A",X"09",X"60",X"2B",X"7E",X"FE",X"FF",
		X"C0",X"06",X"80",X"3A",X"07",X"60",X"FE",X"0B",X"20",X"07",X"3E",X"01",X"32",X"07",X"60",X"18",
		X"15",X"3C",X"F5",X"3A",X"58",X"61",X"FE",X"00",X"28",X"08",X"CD",X"D9",X"0C",X"FE",X"00",X"CA",
		X"19",X"0C",X"F1",X"32",X"07",X"60",X"3A",X"07",X"60",X"FE",X"01",X"C8",X"FE",X"03",X"CC",X"7F",
		X"0E",X"FE",X"05",X"C8",X"FE",X"08",X"CC",X"7F",X"0E",X"FE",X"0A",X"C8",X"FE",X"02",X"CC",X"7F",
		X"0E",X"FE",X"04",X"CC",X"7F",X"0E",X"FE",X"07",X"CC",X"7F",X"0E",X"FE",X"09",X"CC",X"7F",X"0E",
		X"FE",X"06",X"20",X"0C",X"3E",X"12",X"32",X"80",X"65",X"CD",X"7F",X"0E",X"CD",X"60",X"0E",X"C9",
		X"FE",X"0B",X"20",X"0B",X"3E",X"92",X"32",X"80",X"65",X"CD",X"7F",X"0E",X"CD",X"60",X"0E",X"C9",
		X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"27",X"3F",X"CD",X"18",X"20",X"3A",X"58",X"61",
		X"FE",X"00",X"C8",X"3E",X"3F",X"32",X"9C",X"65",X"3A",X"82",X"65",X"32",X"9E",X"65",X"C9",X"F5",
		X"AF",X"32",X"1C",X"60",X"32",X"1D",X"60",X"32",X"1E",X"60",X"78",X"FE",X"80",X"20",X"13",X"3A",
		X"83",X"65",X"3D",X"32",X"83",X"65",X"DD",X"21",X"80",X"65",X"CD",X"72",X"0F",X"CD",X"60",X"0E",
		X"F1",X"C9",X"3A",X"83",X"65",X"3C",X"32",X"83",X"65",X"DD",X"21",X"80",X"65",X"CD",X"72",X"0F",
		X"CD",X"60",X"0E",X"F1",X"C9",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"3A",X"0F",X"91",X"FE",
		X"1E",X"28",X"06",X"3A",X"2F",X"91",X"FE",X"1E",X"C0",X"3A",X"00",X"60",X"FE",X"00",X"C8",X"3A",
		X"54",X"60",X"FE",X"01",X"C8",X"3A",X"26",X"60",X"E6",X"04",X"FE",X"04",X"28",X"1D",X"3A",X"00",
		X"60",X"FE",X"02",X"D8",X"3A",X"51",X"60",X"E6",X"04",X"FE",X"04",X"C0",X"3A",X"00",X"60",X"3D",
		X"27",X"32",X"00",X"60",X"3E",X"02",X"32",X"7D",X"61",X"18",X"05",X"3E",X"01",X"32",X"7D",X"61",
		X"AF",X"32",X"7C",X"61",X"3A",X"00",X"60",X"3D",X"27",X"32",X"00",X"60",X"3E",X"0A",X"32",X"7D",
		X"62",X"32",X"90",X"62",X"CD",X"91",X"35",X"3E",X"01",X"32",X"10",X"62",X"CD",X"94",X"1E",X"CD",
		X"57",X"29",X"3E",X"01",X"32",X"9A",X"60",X"AF",X"32",X"53",X"60",X"32",X"55",X"60",X"3C",X"32",
		X"54",X"60",X"AF",X"21",X"76",X"61",X"06",X"06",X"77",X"23",X"10",X"FC",X"3A",X"63",X"61",X"E6",
		X"03",X"C6",X"01",X"32",X"56",X"60",X"3C",X"32",X"7E",X"61",X"21",X"C2",X"91",X"22",X"C4",X"61",
		X"22",X"FA",X"61",X"3E",X"01",X"32",X"C6",X"61",X"32",X"FC",X"61",X"AF",X"32",X"C7",X"61",X"32",
		X"CF",X"61",X"32",X"14",X"60",X"32",X"1C",X"60",X"32",X"58",X"61",X"CD",X"5B",X"35",X"CD",X"67",
		X"35",X"C9",X"DD",X"7E",X"02",X"D6",X"01",X"E6",X"F8",X"C6",X"04",X"DD",X"77",X"02",X"C9",X"2A",
		X"40",X"61",X"11",X"03",X"00",X"19",X"7E",X"FE",X"FF",X"C8",X"7E",X"47",X"3A",X"42",X"61",X"B8",
		X"C0",X"AF",X"32",X"42",X"61",X"2A",X"40",X"61",X"11",X"25",X"5B",X"CD",X"B2",X"0F",X"3E",X"0F",
		X"D3",X"08",X"3E",X"01",X"32",X"07",X"A0",X"2A",X"40",X"61",X"11",X"04",X"00",X"19",X"22",X"40",
		X"61",X"C9",X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"38",X"D3",X"09",X"0E",X"00",
		X"D5",X"CD",X"CC",X"0F",X"D1",X"EB",X"0E",X"08",X"CD",X"F0",X"0F",X"C9",X"06",X"03",X"79",X"D3",
		X"08",X"7E",X"CD",X"DA",X"0F",X"23",X"0C",X"10",X"F5",X"C9",X"E5",X"87",X"26",X"00",X"6F",X"11",
		X"8F",X"3E",X"19",X"7E",X"D3",X"09",X"0C",X"79",X"D3",X"08",X"23",X"7E",X"D3",X"09",X"E1",X"C9",
		X"06",X"06",X"79",X"D3",X"08",X"0C",X"7E",X"D3",X"09",X"23",X"10",X"F6",X"C9",X"3A",X"43",X"61",
		X"C9",X"06",X"04",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"10",X"F4",X"C9",
		X"3A",X"58",X"61",X"FE",X"00",X"C8",X"3A",X"83",X"65",X"D6",X"02",X"32",X"9F",X"65",X"3A",X"80",
		X"65",X"E6",X"7F",X"FE",X"12",X"C8",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",X"20",X"0E",X"3A",
		X"82",X"65",X"C6",X"08",X"32",X"9E",X"65",X"3E",X"BF",X"32",X"9C",X"65",X"C9",X"3A",X"82",X"65",
		X"D6",X"08",X"32",X"9E",X"65",X"3E",X"3F",X"32",X"9C",X"65",X"C9",X"3A",X"CF",X"61",X"FE",X"00",
		X"C8",X"3A",X"80",X"65",X"E6",X"7F",X"FE",X"1F",X"06",X"37",X"28",X"0D",X"3A",X"80",X"65",X"E6",
		X"7F",X"FE",X"12",X"06",X"37",X"28",X"02",X"06",X"38",X"3A",X"83",X"65",X"32",X"9F",X"65",X"3A",
		X"80",X"65",X"E6",X"7F",X"FE",X"12",X"28",X"16",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",X"28",
		X"0D",X"3A",X"82",X"65",X"C6",X"0C",X"32",X"9E",X"65",X"78",X"32",X"9C",X"65",X"C9",X"3A",X"82",
		X"65",X"D6",X"0C",X"32",X"9E",X"65",X"78",X"F6",X"80",X"32",X"9C",X"65",X"C9",X"3A",X"54",X"60",
		X"FE",X"01",X"28",X"0A",X"3A",X"50",X"60",X"E6",X"80",X"FE",X"80",X"28",X"12",X"C9",X"3A",X"26",
		X"60",X"E6",X"80",X"FE",X"80",X"20",X"0E",X"3A",X"50",X"60",X"E6",X"80",X"FE",X"80",X"C8",X"3E",
		X"01",X"32",X"60",X"61",X"C9",X"3E",X"00",X"32",X"60",X"61",X"C9",X"3E",X"FF",X"FD",X"77",X"03",
		X"C9",X"3A",X"10",X"62",X"FE",X"01",X"C0",X"3A",X"ED",X"61",X"FE",X"01",X"C8",X"3A",X"C0",X"61",
		X"FE",X"01",X"28",X"15",X"21",X"BD",X"61",X"11",X"00",X"A8",X"01",X"06",X"00",X"ED",X"B0",X"AF",
		X"32",X"03",X"A8",X"3E",X"01",X"32",X"C0",X"61",X"C9",X"3E",X"01",X"32",X"03",X"A8",X"C9",X"3A",
		X"C7",X"61",X"FE",X"00",X"C8",X"3A",X"82",X"65",X"C6",X"0E",X"32",X"9E",X"65",X"3A",X"ED",X"61",
		X"FE",X"01",X"28",X"05",X"3E",X"10",X"32",X"9F",X"65",X"3A",X"83",X"65",X"47",X"3A",X"9F",X"65",
		X"B8",X"C8",X"C6",X"01",X"B8",X"C8",X"01",X"C7",X"61",X"D9",X"FD",X"21",X"C4",X"61",X"3E",X"28",
		X"FD",X"77",X"05",X"3E",X"EC",X"FD",X"77",X"06",X"C4",X"BA",X"21",X"C9",X"3A",X"CF",X"61",X"FE",
		X"00",X"C8",X"2A",X"E0",X"61",X"7D",X"FE",X"00",X"20",X"06",X"7C",X"FE",X"00",X"20",X"01",X"C9",
		X"23",X"22",X"E0",X"61",X"11",X"FF",X"01",X"ED",X"52",X"C0",X"21",X"00",X"00",X"22",X"E0",X"61",
		X"3E",X"00",X"DD",X"21",X"CC",X"61",X"DD",X"77",X"03",X"3E",X"FF",X"32",X"9F",X"65",X"C9",X"3A",
		X"99",X"60",X"32",X"98",X"60",X"2A",X"38",X"60",X"22",X"44",X"60",X"FD",X"21",X"57",X"60",X"FD",
		X"22",X"93",X"60",X"DD",X"2A",X"A9",X"04",X"21",X"34",X"60",X"FD",X"21",X"27",X"60",X"CD",X"70",
		X"05",X"3A",X"00",X"B8",X"3A",X"98",X"60",X"32",X"99",X"60",X"C9",X"3A",X"9A",X"60",X"32",X"98",
		X"60",X"2A",X"78",X"60",X"22",X"44",X"60",X"FD",X"21",X"97",X"60",X"FD",X"22",X"93",X"60",X"DD",
		X"2A",X"AB",X"04",X"21",X"74",X"60",X"FD",X"21",X"67",X"60",X"CD",X"70",X"05",X"3A",X"00",X"B8",
		X"3A",X"98",X"60",X"32",X"9A",X"60",X"C9",X"BF",X"73",X"FB",X"EE",X"8B",X"B8",X"AF",X"BB",X"7C",
		X"52",X"9B",X"FC",X"BF",X"7D",X"B6",X"E3",X"5F",X"EE",X"BB",X"FB",X"7B",X"0F",X"AE",X"F9",X"FE",
		X"95",X"BB",X"FF",X"BF",X"13",X"BF",X"FF",X"9A",X"BB",X"BE",X"9F",X"B5",X"EA",X"3E",X"ED",X"DF",
		X"67",X"EB",X"BB",X"BC",X"1C",X"CF",X"7A",X"36",X"D3",X"6E",X"20",X"FF",X"74",X"BF",X"97",X"7E",
		X"AF",X"32",X"00",X"A0",X"F3",X"3C",X"C3",X"80",X"24",X"21",X"00",X"05",X"CD",X"38",X"2C",X"3E",
		X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3E",X"40",X"32",X"E8",X"61",X"CD",X"00",X"37",X"CD",
		X"5B",X"35",X"CD",X"67",X"35",X"21",X"3C",X"51",X"22",X"40",X"61",X"F3",X"3A",X"00",X"B8",X"CD",
		X"94",X"1E",X"CD",X"57",X"29",X"AF",X"32",X"25",X"60",X"3C",X"32",X"9A",X"60",X"3E",X"03",X"32",
		X"99",X"60",X"3E",X"01",X"ED",X"56",X"32",X"00",X"A0",X"FB",X"3A",X"00",X"A8",X"CD",X"CF",X"34",
		X"CD",X"A4",X"24",X"DD",X"21",X"80",X"65",X"FD",X"21",X"94",X"65",X"11",X"04",X"00",X"3A",X"0D",
		X"60",X"47",X"3A",X"99",X"60",X"B8",X"20",X"13",X"CD",X"37",X"55",X"FE",X"00",X"28",X"0C",X"3A",
		X"56",X"61",X"FE",X"00",X"20",X"05",X"3E",X"01",X"32",X"25",X"60",X"DD",X"21",X"80",X"65",X"FD",
		X"21",X"98",X"65",X"11",X"04",X"00",X"CD",X"53",X"16",X"3A",X"0D",X"60",X"47",X"3A",X"9A",X"60",
		X"B8",X"20",X"13",X"CD",X"37",X"55",X"FE",X"00",X"28",X"0C",X"3A",X"57",X"61",X"FE",X"00",X"20",
		X"05",X"3E",X"01",X"32",X"25",X"60",X"3A",X"54",X"60",X"FE",X"01",X"28",X"63",X"3E",X"01",X"32",
		X"01",X"A0",X"32",X"02",X"A0",X"3A",X"53",X"60",X"FE",X"01",X"20",X"54",X"3A",X"10",X"62",X"FE",
		X"01",X"28",X"4D",X"F3",X"3A",X"55",X"60",X"FE",X"01",X"28",X"1F",X"3A",X"00",X"B8",X"CD",X"2C",
		X"2A",X"CD",X"EC",X"1D",X"CD",X"BE",X"39",X"21",X"3C",X"51",X"22",X"40",X"61",X"3E",X"01",X"32",
		X"55",X"60",X"3A",X"54",X"60",X"FE",X"01",X"CA",X"42",X"12",X"3A",X"10",X"62",X"FE",X"01",X"28",
		X"1F",X"3A",X"00",X"60",X"FE",X"01",X"20",X"0C",X"11",X"DF",X"56",X"21",X"11",X"93",X"CD",X"F9",
		X"30",X"C3",X"42",X"12",X"11",X"F2",X"56",X"21",X"11",X"93",X"CD",X"F9",X"30",X"C3",X"42",X"12",
		X"CD",X"3F",X"1E",X"FE",X"01",X"CA",X"2B",X"12",X"3A",X"E8",X"61",X"FE",X"00",X"20",X"08",X"CD",
		X"70",X"1E",X"FE",X"01",X"CA",X"2B",X"12",X"CD",X"7A",X"1E",X"32",X"00",X"B8",X"CD",X"30",X"1C",
		X"3A",X"A3",X"58",X"32",X"73",X"62",X"3A",X"00",X"B8",X"3A",X"0D",X"60",X"47",X"3A",X"99",X"60",
		X"B8",X"CC",X"38",X"1B",X"FB",X"CD",X"C9",X"1C",X"3A",X"0F",X"57",X"32",X"70",X"62",X"3A",X"00",
		X"B8",X"3A",X"00",X"B8",X"3A",X"0D",X"60",X"47",X"3A",X"9A",X"60",X"B8",X"CC",X"94",X"1C",X"FB",
		X"CD",X"B3",X"25",X"32",X"00",X"B0",X"3A",X"99",X"60",X"32",X"98",X"60",X"FD",X"21",X"94",X"65",
		X"FD",X"22",X"93",X"60",X"DD",X"21",X"27",X"60",X"DD",X"22",X"95",X"60",X"DD",X"21",X"35",X"60",
		X"FD",X"21",X"94",X"65",X"ED",X"5B",X"38",X"60",X"ED",X"53",X"91",X"60",X"3A",X"00",X"B8",X"CD",
		X"D1",X"19",X"DD",X"21",X"3B",X"60",X"21",X"57",X"60",X"11",X"48",X"61",X"CD",X"08",X"19",X"3A",
		X"48",X"61",X"FE",X"00",X"20",X"2D",X"3A",X"57",X"60",X"FE",X"F0",X"D4",X"A3",X"31",X"FE",X"10",
		X"FD",X"21",X"94",X"65",X"FD",X"22",X"93",X"60",X"DD",X"21",X"27",X"60",X"DD",X"22",X"95",X"60",
		X"FD",X"21",X"94",X"65",X"ED",X"5B",X"38",X"60",X"ED",X"53",X"91",X"60",X"DD",X"21",X"35",X"60",
		X"D4",X"23",X"21",X"3A",X"9A",X"60",X"32",X"98",X"60",X"FD",X"21",X"98",X"65",X"FD",X"22",X"93",
		X"60",X"DD",X"21",X"67",X"60",X"DD",X"22",X"95",X"60",X"DD",X"21",X"75",X"60",X"FD",X"21",X"98",
		X"65",X"ED",X"5B",X"78",X"60",X"ED",X"53",X"91",X"60",X"3A",X"00",X"B8",X"3A",X"0C",X"57",X"32",
		X"71",X"62",X"CD",X"D1",X"19",X"DD",X"21",X"7B",X"60",X"21",X"97",X"60",X"11",X"49",X"61",X"CD",
		X"08",X"19",X"CD",X"53",X"16",X"3A",X"49",X"61",X"FE",X"00",X"20",X"2D",X"3A",X"97",X"60",X"FE",
		X"F0",X"D4",X"C1",X"31",X"FE",X"10",X"FD",X"21",X"98",X"65",X"FD",X"22",X"93",X"60",X"DD",X"21",
		X"67",X"60",X"DD",X"22",X"95",X"60",X"FD",X"21",X"98",X"65",X"ED",X"5B",X"78",X"60",X"ED",X"53",
		X"91",X"60",X"DD",X"21",X"75",X"60",X"D4",X"23",X"21",X"FB",X"CD",X"75",X"55",X"7E",X"FE",X"E0",
		X"CA",X"55",X"14",X"18",X"05",X"3E",X"01",X"32",X"77",X"60",X"CD",X"68",X"55",X"7E",X"FE",X"E0",
		X"28",X"02",X"18",X"05",X"3E",X"01",X"32",X"37",X"60",X"2A",X"38",X"60",X"FD",X"21",X"37",X"60",
		X"DD",X"21",X"94",X"65",X"CD",X"05",X"26",X"2A",X"38",X"60",X"DD",X"21",X"94",X"65",X"CD",X"0E",
		X"25",X"2A",X"78",X"60",X"FD",X"21",X"77",X"60",X"DD",X"21",X"98",X"65",X"CD",X"05",X"26",X"2A",
		X"78",X"60",X"DD",X"21",X"98",X"65",X"CD",X"0E",X"25",X"3A",X"00",X"B8",X"CD",X"5E",X"55",X"FB",
		X"7E",X"FE",X"E0",X"28",X"0E",X"3A",X"4E",X"60",X"FE",X"01",X"28",X"0C",X"3E",X"00",X"32",X"08",
		X"60",X"18",X"05",X"3E",X"01",X"32",X"08",X"60",X"2A",X"09",X"60",X"FD",X"21",X"08",X"60",X"DD",
		X"21",X"80",X"65",X"CD",X"05",X"26",X"2A",X"09",X"60",X"DD",X"21",X"80",X"65",X"CD",X"0E",X"25",
		X"3E",X"01",X"32",X"6F",X"62",X"3A",X"00",X"B8",X"CD",X"28",X"2C",X"CD",X"19",X"32",X"3E",X"00",
		X"32",X"6F",X"62",X"CD",X"84",X"1D",X"CD",X"73",X"1D",X"FE",X"01",X"CA",X"2B",X"12",X"DD",X"21",
		X"3C",X"60",X"06",X"04",X"DD",X"7E",X"00",X"FE",X"00",X"20",X"2A",X"DD",X"23",X"10",X"F5",X"21",
		X"27",X"60",X"22",X"95",X"60",X"21",X"44",X"61",X"22",X"46",X"61",X"3A",X"99",X"60",X"32",X"98",
		X"60",X"DD",X"21",X"80",X"65",X"FD",X"21",X"94",X"65",X"ED",X"5B",X"38",X"60",X"21",X"3B",X"60",
		X"CD",X"FA",X"2A",X"18",X"04",X"AF",X"32",X"48",X"61",X"DD",X"21",X"7C",X"60",X"06",X"04",X"DD",
		X"7E",X"00",X"FE",X"00",X"20",X"2A",X"DD",X"23",X"10",X"F5",X"21",X"67",X"60",X"22",X"95",X"60",
		X"21",X"45",X"61",X"22",X"46",X"61",X"3A",X"9A",X"60",X"32",X"98",X"60",X"DD",X"21",X"80",X"65",
		X"FD",X"21",X"98",X"65",X"ED",X"5B",X"78",X"60",X"21",X"7B",X"60",X"CD",X"FA",X"2A",X"18",X"04",
		X"AF",X"32",X"49",X"61",X"FB",X"CD",X"DE",X"17",X"CD",X"53",X"16",X"3A",X"CF",X"61",X"FE",X"01",
		X"28",X"21",X"3A",X"58",X"61",X"FE",X"01",X"28",X"1A",X"01",X"C7",X"61",X"FD",X"21",X"C4",X"61",
		X"3E",X"3A",X"FD",X"77",X"04",X"3E",X"28",X"FD",X"77",X"05",X"3E",X"EC",X"32",X"CA",X"61",X"F3",
		X"CD",X"37",X"21",X"F3",X"06",X"04",X"FD",X"21",X"D0",X"61",X"3A",X"C7",X"61",X"FE",X"01",X"CA",
		X"CF",X"15",X"C5",X"FD",X"E5",X"01",X"CF",X"61",X"FD",X"21",X"CC",X"61",X"3E",X"37",X"FD",X"77",
		X"04",X"3E",X"20",X"FD",X"77",X"05",X"3A",X"00",X"B8",X"3E",X"E4",X"32",X"D2",X"61",X"CD",X"37",
		X"21",X"FD",X"E1",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"CD",X"B7",X"22",X"C1",X"10",X"D3",X"FB",
		X"3A",X"CF",X"61",X"FE",X"00",X"28",X"4A",X"3A",X"99",X"60",X"47",X"3A",X"70",X"62",X"B8",X"3A",
		X"0D",X"60",X"B8",X"20",X"19",X"DD",X"21",X"94",X"65",X"FD",X"21",X"9C",X"65",X"0E",X"00",X"06",
		X"06",X"CD",X"D5",X"2A",X"FE",X"01",X"20",X"06",X"CD",X"41",X"22",X"CD",X"3D",X"31",X"DD",X"21",
		X"98",X"65",X"FD",X"21",X"9C",X"65",X"3A",X"9A",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"20",X"11",
		X"0E",X"00",X"06",X"06",X"CD",X"D5",X"2A",X"FE",X"01",X"20",X"06",X"CD",X"7C",X"22",X"CD",X"3D",
		X"31",X"DD",X"21",X"80",X"65",X"FD",X"21",X"84",X"65",X"CD",X"D1",X"2A",X"FE",X"01",X"20",X"11",
		X"3E",X"01",X"32",X"25",X"60",X"AF",X"32",X"29",X"60",X"CD",X"73",X"1D",X"FE",X"01",X"CA",X"2B",
		X"12",X"FB",X"CD",X"4D",X"2C",X"CD",X"A1",X"3B",X"3A",X"ED",X"61",X"FE",X"00",X"CC",X"DC",X"22",
		X"C3",X"42",X"12",X"3A",X"ED",X"61",X"FE",X"00",X"C0",X"3A",X"7F",X"62",X"FE",X"01",X"C0",X"E5",
		X"D5",X"F5",X"C5",X"FD",X"E5",X"DD",X"E5",X"3A",X"98",X"60",X"32",X"80",X"62",X"CD",X"BC",X"3B",
		X"AF",X"32",X"7F",X"62",X"3A",X"80",X"62",X"32",X"98",X"60",X"DD",X"E1",X"FD",X"E1",X"C1",X"F1",
		X"D1",X"E1",X"C9",X"3A",X"5E",X"61",X"FE",X"00",X"20",X"06",X"3A",X"59",X"61",X"FE",X"00",X"C8",
		X"DD",X"21",X"9C",X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",X"32",X"98",X"60",X"DD",X"35",
		X"03",X"CD",X"8C",X"55",X"FB",X"DD",X"21",X"9C",X"65",X"DD",X"34",X"03",X"FB",X"7E",X"E5",X"21",
		X"24",X"5B",X"01",X"07",X"00",X"ED",X"B9",X"E1",X"C2",X"C5",X"16",X"3E",X"01",X"32",X"5E",X"61",
		X"AF",X"32",X"59",X"61",X"C9",X"AF",X"32",X"5E",X"61",X"3C",X"32",X"59",X"61",X"DD",X"21",X"9C",
		X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",X"8C",X"55",X"FB",X"7E",
		X"E5",X"21",X"D0",X"17",X"01",X"22",X"00",X"ED",X"B9",X"E1",X"C8",X"AF",X"32",X"5E",X"61",X"32",
		X"59",X"61",X"FD",X"2A",X"5C",X"61",X"3A",X"0D",X"60",X"FD",X"77",X"02",X"FE",X"01",X"20",X"05",
		X"7C",X"C6",X"50",X"18",X"0C",X"FE",X"02",X"20",X"05",X"7C",X"C6",X"4C",X"18",X"03",X"7C",X"C6",
		X"48",X"67",X"AF",X"7D",X"D6",X"22",X"6F",X"7C",X"DE",X"00",X"67",X"7E",X"FE",X"D0",X"28",X"10",
		X"EB",X"21",X"D0",X"17",X"01",X"07",X"00",X"ED",X"B9",X"EB",X"28",X"04",X"11",X"20",X"00",X"19",
		X"F3",X"FD",X"75",X"00",X"7D",X"FE",X"C0",X"20",X"02",X"3E",X"68",X"FD",X"74",X"01",X"3A",X"0D",
		X"60",X"FD",X"77",X"02",X"FB",X"23",X"7E",X"FE",X"ED",X"28",X"13",X"FE",X"EF",X"28",X"0F",X"7D",
		X"C6",X"20",X"6F",X"7C",X"CE",X"00",X"67",X"7E",X"FE",X"ED",X"28",X"02",X"18",X"42",X"DD",X"E5",
		X"CD",X"D5",X"17",X"3A",X"9D",X"65",X"FE",X"24",X"20",X"0B",X"3E",X"20",X"32",X"9D",X"65",X"CD",
		X"D5",X"17",X"CD",X"D5",X"17",X"21",X"1B",X"3F",X"CD",X"18",X"20",X"CD",X"EB",X"3D",X"20",X"0A",
		X"21",X"78",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"DD",X"E1",X"F3",X"AF",X"FD",X"77",
		X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FB",X"3E",X"40",X"32",X"E8",X"61",X"CD",X"00",X"3B",
		X"AF",X"DD",X"21",X"9C",X"65",X"DD",X"77",X"02",X"3E",X"FF",X"DD",X"77",X"03",X"C9",X"49",X"FA",
		X"FD",X"7E",X"67",X"98",X"FC",X"BA",X"CF",X"74",X"6F",X"6D",X"6B",X"87",X"E5",X"E0",X"9B",X"FD",
		X"70",X"3D",X"41",X"63",X"1B",X"1A",X"27",X"26",X"25",X"24",X"FF",X"DF",X"E0",X"4A",X"DE",X"4B",
		X"DE",X"E2",X"C2",X"A2",X"E2",X"2A",X"E7",X"61",X"2E",X"00",X"CD",X"90",X"5C",X"C9",X"3A",X"58",
		X"61",X"FE",X"00",X"C2",X"5F",X"19",X"3A",X"CF",X"61",X"FE",X"01",X"C8",X"3A",X"C7",X"61",X"FE",
		X"01",X"C8",X"3A",X"59",X"61",X"FE",X"01",X"C8",X"3A",X"5E",X"61",X"FE",X"01",X"C8",X"FD",X"21",
		X"9C",X"60",X"06",X"12",X"2A",X"09",X"60",X"3E",X"24",X"32",X"7B",X"62",X"FD",X"7E",X"02",X"C5",
		X"47",X"3A",X"0D",X"60",X"B8",X"C1",X"C2",X"30",X"18",X"FD",X"56",X"01",X"FD",X"5E",X"00",X"13",
		X"13",X"CD",X"45",X"19",X"AF",X"E5",X"ED",X"52",X"E1",X"28",X"13",X"CD",X"85",X"35",X"28",X"0E",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"3E",X"20",X"32",X"7B",X"62",X"10",X"CF",X"C9",X"CD",X"A4",
		X"19",X"78",X"FE",X"00",X"C8",X"3A",X"CF",X"61",X"FE",X"00",X"28",X"1F",X"FD",X"E5",X"E5",X"01",
		X"CF",X"61",X"FD",X"21",X"CC",X"61",X"3E",X"38",X"FD",X"77",X"04",X"3E",X"28",X"FD",X"77",X"05",
		X"3E",X"E4",X"32",X"D2",X"61",X"CD",X"BA",X"21",X"E1",X"FD",X"E1",X"DD",X"21",X"80",X"65",X"3E",
		X"3F",X"DD",X"77",X"1C",X"3A",X"7B",X"62",X"DD",X"77",X"1D",X"DD",X"7E",X"03",X"DD",X"77",X"1F",
		X"DD",X"7E",X"02",X"D6",X"08",X"DD",X"77",X"1E",X"CD",X"EB",X"3D",X"20",X"0A",X"21",X"A8",X"5B",
		X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"3E",X"01",X"32",X"58",X"61",X"FD",X"22",X"5C",X"61",
		X"FD",X"66",X"01",X"FD",X"6E",X"00",X"22",X"F6",X"61",X"AF",X"32",X"7E",X"62",X"F3",X"FD",X"77",
		X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FB",X"3A",X"7B",X"62",X"FE",X"24",X"3E",X"00",X"20",
		X"02",X"3E",X"01",X"32",X"7C",X"62",X"C9",X"3A",X"7E",X"62",X"FE",X"07",X"D0",X"2A",X"F6",X"61",
		X"7C",X"FE",X"00",X"C8",X"7D",X"E6",X"0F",X"FE",X"00",X"C8",X"CD",X"2F",X"19",X"CD",X"15",X"19",
		X"23",X"CD",X"2F",X"19",X"CD",X"15",X"19",X"11",X"20",X"00",X"19",X"CD",X"2F",X"19",X"CD",X"15",
		X"19",X"2B",X"CD",X"2F",X"19",X"CD",X"15",X"19",X"3A",X"7E",X"62",X"3C",X"32",X"7E",X"62",X"3A",
		X"0D",X"60",X"FE",X"02",X"CC",X"E3",X"33",X"C9",X"DD",X"7E",X"00",X"FE",X"01",X"C8",X"7E",X"FE",
		X"F0",X"D8",X"AF",X"12",X"C9",X"06",X"1F",X"7E",X"FE",X"49",X"28",X"0A",X"FE",X"4A",X"28",X"06",
		X"FE",X"4B",X"28",X"02",X"06",X"3F",X"E5",X"7C",X"C6",X"08",X"67",X"78",X"77",X"E1",X"C9",X"7C",
		X"57",X"7D",X"5F",X"CD",X"45",X"19",X"1A",X"77",X"1A",X"BE",X"20",X"FA",X"E5",X"7C",X"C6",X"08",
		X"67",X"AF",X"77",X"E1",X"C9",X"3A",X"0D",X"60",X"FE",X"01",X"20",X"05",X"7A",X"D6",X"50",X"57",
		X"C9",X"FE",X"02",X"20",X"05",X"7A",X"D6",X"4C",X"57",X"C9",X"7A",X"D6",X"48",X"57",X"C9",X"3A",
		X"9E",X"65",X"FE",X"E0",X"D0",X"FE",X"18",X"D8",X"CD",X"A4",X"19",X"78",X"FE",X"00",X"C8",X"DD",
		X"21",X"9C",X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",X"8C",X"55",
		X"FB",X"2B",X"7E",X"E5",X"CD",X"B3",X"19",X"E1",X"C0",X"2B",X"E5",X"CD",X"B3",X"19",X"E1",X"C0",
		X"11",X"21",X"00",X"19",X"CD",X"B3",X"19",X"C0",X"AF",X"32",X"58",X"61",X"32",X"7C",X"62",X"3C",
		X"32",X"59",X"61",X"C9",X"06",X"00",X"3A",X"60",X"61",X"FE",X"00",X"C8",X"AF",X"32",X"60",X"61",
		X"06",X"01",X"C9",X"21",X"D0",X"19",X"01",X"15",X"00",X"ED",X"B9",X"C9",X"FF",X"F0",X"F1",X"F2",
		X"F3",X"F4",X"F5",X"F6",X"F7",X"EF",X"EE",X"ED",X"EC",X"EB",X"EA",X"DF",X"DE",X"4A",X"49",X"4B",
		X"E0",X"FD",X"E5",X"FD",X"21",X"74",X"59",X"FD",X"7E",X"00",X"67",X"FD",X"7E",X"01",X"6F",X"AF",
		X"ED",X"52",X"28",X"17",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"3A",X"00",X"B8",X"FD",X"7E",X"02",
		X"FE",X"FF",X"20",X"E3",X"AF",X"DD",X"77",X"11",X"FD",X"E1",X"C9",X"DD",X"E5",X"FD",X"22",X"4B",
		X"60",X"3A",X"98",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"28",X"03",X"CD",X"BD",X"1B",X"06",X"08",
		X"DD",X"7E",X"11",X"FE",X"01",X"CA",X"0B",X"1B",X"DD",X"7E",X"07",X"FE",X"00",X"C2",X"0B",X"1B",
		X"DD",X"23",X"10",X"F4",X"DD",X"E1",X"AF",X"DD",X"77",X"15",X"3A",X"47",X"60",X"FE",X"00",X"CA",
		X"5C",X"1A",X"3A",X"82",X"65",X"47",X"FD",X"E1",X"FD",X"7E",X"02",X"FD",X"E5",X"B8",X"F5",X"D4",
		X"10",X"1B",X"F1",X"DC",X"19",X"1B",X"3A",X"83",X"65",X"47",X"FD",X"E1",X"FD",X"7E",X"03",X"FD",
		X"E5",X"B8",X"F5",X"DC",X"2B",X"1B",X"F1",X"D4",X"22",X"1B",X"18",X"58",X"3A",X"00",X"A0",X"E5",
		X"21",X"34",X"1B",X"E6",X"03",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"3A",X"00",X"B8",X"7E",X"C5",
		X"DD",X"E5",X"DD",X"2A",X"95",X"60",X"47",X"DD",X"7E",X"00",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",
		X"CB",X"0F",X"E6",X"0F",X"FE",X"01",X"20",X"04",X"3E",X"02",X"18",X"16",X"FE",X"02",X"20",X"04",
		X"3E",X"01",X"18",X"0E",X"FE",X"04",X"20",X"04",X"3E",X"08",X"18",X"06",X"FE",X"08",X"20",X"02",
		X"3E",X"04",X"B8",X"20",X"07",X"DD",X"E1",X"C1",X"E1",X"C3",X"5C",X"1A",X"DD",X"E1",X"78",X"C1",
		X"E1",X"DD",X"77",X"15",X"AF",X"FD",X"2A",X"4B",X"60",X"FD",X"7E",X"02",X"CB",X"0F",X"CB",X"0F",
		X"CB",X"0F",X"CB",X"0F",X"47",X"DD",X"7E",X"15",X"A0",X"CB",X"0F",X"2A",X"91",X"60",X"32",X"44",
		X"60",X"FD",X"21",X"94",X"65",X"FD",X"22",X"93",X"60",X"2A",X"95",X"60",X"30",X"05",X"CD",X"B3",
		X"1B",X"18",X"20",X"CB",X"0F",X"30",X"05",X"CD",X"A9",X"1B",X"18",X"17",X"CB",X"0F",X"30",X"05",
		X"CD",X"8B",X"1B",X"18",X"07",X"CB",X"0F",X"30",X"0A",X"CD",X"6D",X"1B",X"3A",X"0B",X"60",X"FE",
		X"02",X"20",X"05",X"3E",X"01",X"DD",X"77",X"11",X"FD",X"E1",X"C9",X"DD",X"E1",X"FD",X"E1",X"C9",
		X"DD",X"7E",X"15",X"F6",X"04",X"DD",X"77",X"15",X"C9",X"DD",X"7E",X"15",X"F6",X"08",X"DD",X"77",
		X"15",X"C9",X"DD",X"7E",X"15",X"F6",X"01",X"DD",X"77",X"15",X"C9",X"DD",X"7E",X"15",X"F6",X"02",
		X"DD",X"77",X"15",X"C9",X"08",X"04",X"02",X"01",X"2A",X"38",X"60",X"22",X"91",X"60",X"FD",X"21",
		X"94",X"65",X"FD",X"22",X"93",X"60",X"21",X"27",X"60",X"22",X"95",X"60",X"3A",X"3C",X"60",X"FE",
		X"00",X"C4",X"6D",X"1B",X"3A",X"3D",X"60",X"FE",X"00",X"C4",X"8B",X"1B",X"3A",X"3E",X"60",X"FE",
		X"00",X"C4",X"B3",X"1B",X"3A",X"3F",X"60",X"FE",X"00",X"C4",X"A9",X"1B",X"C9",X"2A",X"91",X"60",
		X"DD",X"E5",X"DD",X"2A",X"93",X"60",X"CD",X"FA",X"0C",X"DD",X"E1",X"3A",X"0B",X"60",X"FE",X"02",
		X"C0",X"E5",X"2A",X"95",X"60",X"AF",X"CB",X"FF",X"77",X"E1",X"C9",X"2A",X"91",X"60",X"DD",X"E5",
		X"DD",X"2A",X"93",X"60",X"CD",X"69",X"0D",X"DD",X"E1",X"3A",X"0B",X"60",X"FE",X"02",X"C0",X"E5",
		X"2A",X"95",X"60",X"AF",X"CB",X"F7",X"77",X"E1",X"C9",X"AF",X"E5",X"2A",X"95",X"60",X"CB",X"EF",
		X"77",X"E1",X"C9",X"AF",X"E5",X"2A",X"95",X"60",X"CB",X"E7",X"77",X"E1",X"C9",X"DD",X"E5",X"FD",
		X"E5",X"E5",X"C5",X"D5",X"78",X"FE",X"01",X"20",X"06",X"FD",X"21",X"10",X"5A",X"18",X"1B",X"FE",
		X"02",X"20",X"13",X"47",X"3A",X"0D",X"60",X"B8",X"30",X"06",X"FD",X"21",X"3D",X"5A",X"18",X"0A",
		X"FD",X"21",X"76",X"5A",X"18",X"04",X"FD",X"21",X"AF",X"5A",X"D1",X"FD",X"7E",X"00",X"67",X"FD",
		X"7E",X"01",X"6F",X"AF",X"ED",X"52",X"28",X"10",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"7E",
		X"02",X"FE",X"FF",X"20",X"E6",X"C3",X"26",X"1C",X"FD",X"7E",X"02",X"FE",X"80",X"20",X"06",X"CD",
		X"6D",X"1B",X"C3",X"26",X"1C",X"FE",X"40",X"20",X"06",X"CD",X"8B",X"1B",X"C3",X"26",X"1C",X"DD",
		X"2A",X"95",X"60",X"DD",X"77",X"00",X"C1",X"E1",X"FD",X"E1",X"DD",X"E1",X"E1",X"C3",X"0B",X"1B",
		X"3A",X"0D",X"60",X"47",X"3A",X"99",X"60",X"B8",X"C0",X"DD",X"21",X"3D",X"60",X"2A",X"38",X"60",
		X"01",X"E0",X"FF",X"3A",X"CF",X"61",X"FE",X"00",X"3E",X"40",X"20",X"06",X"DD",X"21",X"3C",X"60",
		X"3E",X"80",X"08",X"CD",X"33",X"1D",X"2A",X"38",X"60",X"DD",X"21",X"3C",X"60",X"01",X"20",X"00",
		X"3A",X"CF",X"61",X"FE",X"00",X"3E",X"80",X"20",X"06",X"DD",X"21",X"3D",X"60",X"3E",X"40",X"08",
		X"CD",X"33",X"1D",X"2A",X"38",X"60",X"01",X"FF",X"FF",X"3E",X"10",X"08",X"DD",X"21",X"3E",X"60",
		X"CD",X"33",X"1D",X"2A",X"38",X"60",X"DD",X"21",X"3F",X"60",X"01",X"01",X"00",X"3E",X"20",X"08",
		X"CD",X"33",X"1D",X"C9",X"2A",X"78",X"60",X"22",X"91",X"60",X"FD",X"21",X"98",X"65",X"FD",X"22",
		X"93",X"60",X"21",X"67",X"60",X"22",X"95",X"60",X"3A",X"7C",X"60",X"FE",X"00",X"C4",X"6D",X"1B",
		X"3A",X"7D",X"60",X"FE",X"00",X"C4",X"8B",X"1B",X"3A",X"7E",X"60",X"FE",X"00",X"C4",X"B3",X"1B",
		X"3A",X"7F",X"60",X"FE",X"00",X"C4",X"A9",X"1B",X"C9",X"3A",X"0D",X"60",X"47",X"3A",X"9A",X"60",
		X"B8",X"C0",X"DD",X"21",X"7D",X"60",X"2A",X"78",X"60",X"01",X"E0",X"FF",X"3A",X"CF",X"61",X"FE",
		X"00",X"3E",X"40",X"20",X"06",X"DD",X"21",X"7C",X"60",X"3E",X"80",X"08",X"CD",X"33",X"1D",X"2A",
		X"78",X"60",X"01",X"20",X"00",X"DD",X"21",X"7C",X"60",X"3A",X"CF",X"61",X"FE",X"00",X"3A",X"B2",
		X"91",X"32",X"72",X"62",X"3E",X"80",X"20",X"06",X"DD",X"21",X"7D",X"60",X"3E",X"40",X"08",X"CD",
		X"33",X"1D",X"2A",X"78",X"60",X"01",X"FF",X"FF",X"3E",X"10",X"08",X"DD",X"21",X"7E",X"60",X"CD",
		X"33",X"1D",X"2A",X"78",X"60",X"DD",X"21",X"7F",X"60",X"01",X"01",X"00",X"3E",X"20",X"08",X"CD",
		X"33",X"1D",X"C9",X"2B",X"2B",X"AF",X"DD",X"77",X"00",X"ED",X"4A",X"7E",X"C5",X"06",X"08",X"FD",
		X"21",X"6B",X"1D",X"FD",X"BE",X"00",X"28",X"06",X"FD",X"23",X"10",X"F7",X"C1",X"C9",X"C1",X"E5",
		X"ED",X"5B",X"09",X"60",X"1B",X"1B",X"AF",X"ED",X"52",X"E1",X"28",X"0A",X"E5",X"13",X"AF",X"ED",
		X"52",X"E1",X"28",X"02",X"18",X"CF",X"08",X"DD",X"77",X"00",X"C9",X"E0",X"FF",X"DF",X"DE",X"DE",
		X"49",X"4A",X"4B",X"3A",X"29",X"60",X"FE",X"01",X"28",X"08",X"3A",X"25",X"60",X"FE",X"01",X"CA",
		X"50",X"1F",X"AF",X"C9",X"3A",X"25",X"60",X"FE",X"01",X"C8",X"3A",X"29",X"60",X"FE",X"01",X"C8",
		X"DD",X"21",X"82",X"65",X"FD",X"21",X"8A",X"65",X"21",X"22",X"60",X"11",X"04",X"00",X"3A",X"2A",
		X"60",X"FE",X"01",X"C8",X"CD",X"B4",X"1D",X"23",X"FD",X"19",X"CD",X"B4",X"1D",X"23",X"FD",X"19",
		X"CD",X"B4",X"1D",X"C9",X"DD",X"7E",X"01",X"3C",X"FD",X"BE",X"01",X"C0",X"FD",X"7E",X"00",X"D6",
		X"0D",X"47",X"C6",X"04",X"4F",X"CD",X"DE",X"1D",X"32",X"25",X"60",X"FE",X"01",X"C8",X"FD",X"7E",
		X"00",X"C6",X"0A",X"47",X"C6",X"04",X"4F",X"CD",X"DE",X"1D",X"32",X"25",X"60",X"C9",X"DD",X"7E",
		X"00",X"B8",X"38",X"06",X"B9",X"30",X"03",X"3E",X"01",X"C9",X"AF",X"C9",X"11",X"80",X"56",X"21",
		X"A0",X"93",X"CD",X"F9",X"30",X"11",X"80",X"56",X"21",X"20",X"91",X"CD",X"F9",X"30",X"11",X"05",
		X"57",X"21",X"40",X"92",X"CD",X"F9",X"30",X"3E",X"02",X"21",X"40",X"90",X"77",X"11",X"89",X"56",
		X"21",X"9F",X"91",X"CD",X"F9",X"30",X"3A",X"04",X"60",X"32",X"9F",X"90",X"3A",X"05",X"60",X"32",
		X"BF",X"90",X"CD",X"26",X"1E",X"C9",X"3E",X"02",X"21",X"40",X"98",X"CD",X"05",X"56",X"3E",X"08",
		X"21",X"5F",X"98",X"CD",X"05",X"56",X"3E",X"05",X"21",X"41",X"98",X"CD",X"05",X"56",X"C9",X"3A",
		X"4D",X"60",X"FE",X"12",X"38",X"1E",X"3E",X"01",X"32",X"4E",X"60",X"2A",X"09",X"60",X"7E",X"FE",
		X"F8",X"E5",X"21",X"67",X"1E",X"01",X"02",X"00",X"ED",X"B9",X"E1",X"20",X"0B",X"3A",X"14",X"60",
		X"FE",X"01",X"28",X"0C",X"AF",X"C9",X"FB",X"E0",X"3A",X"83",X"65",X"D6",X"02",X"32",X"83",X"65",
		X"AF",X"32",X"08",X"60",X"CD",X"50",X"1F",X"3E",X"01",X"C9",X"3A",X"54",X"60",X"FE",X"01",X"28",
		X"0C",X"3A",X"00",X"60",X"FE",X"00",X"28",X"06",X"3E",X"01",X"32",X"53",X"60",X"C9",X"3E",X"00",
		X"32",X"53",X"60",X"C9",X"3A",X"10",X"62",X"FE",X"01",X"20",X"0F",X"CD",X"EB",X"3D",X"20",X"0A",
		X"21",X"00",X"50",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"AF",X"32",X"03",X"A0",X"CD",X"4C",
		X"28",X"3E",X"01",X"32",X"16",X"60",X"CD",X"EC",X"1D",X"3E",X"01",X"32",X"0D",X"60",X"32",X"03",
		X"A0",X"3E",X"20",X"21",X"80",X"65",X"77",X"23",X"3E",X"08",X"77",X"23",X"3E",X"29",X"77",X"23",
		X"3E",X"E0",X"77",X"32",X"29",X"60",X"3E",X"40",X"32",X"65",X"61",X"3E",X"C8",X"32",X"66",X"61",
		X"11",X"C7",X"61",X"21",X"38",X"1F",X"01",X"18",X"00",X"ED",X"B0",X"3E",X"40",X"32",X"E8",X"61",
		X"3E",X"01",X"32",X"86",X"62",X"32",X"19",X"60",X"3E",X"B0",X"32",X"9A",X"65",X"AF",X"32",X"97",
		X"60",X"32",X"88",X"62",X"32",X"08",X"60",X"32",X"13",X"60",X"32",X"29",X"60",X"32",X"2A",X"60",
		X"32",X"4E",X"60",X"32",X"77",X"60",X"32",X"28",X"60",X"32",X"E0",X"61",X"32",X"E1",X"61",X"32",
		X"14",X"60",X"32",X"13",X"60",X"3A",X"C4",X"61",X"FE",X"00",X"28",X"05",X"E6",X"02",X"FE",X"02",
		X"C8",X"21",X"C2",X"91",X"22",X"C4",X"61",X"C9",X"00",X"00",X"00",X"00",X"00",X"55",X"92",X"03",
		X"00",X"00",X"00",X"00",X"58",X"91",X"01",X"D1",X"92",X"02",X"28",X"91",X"01",X"A2",X"90",X"02",
		X"3E",X"01",X"32",X"F1",X"61",X"CD",X"8C",X"3B",X"79",X"FE",X"01",X"CC",X"4F",X"35",X"3A",X"7C",
		X"61",X"32",X"6C",X"62",X"2A",X"09",X"60",X"FD",X"21",X"08",X"60",X"DD",X"21",X"80",X"65",X"CD",
		X"05",X"26",X"3E",X"01",X"32",X"51",X"61",X"32",X"00",X"A0",X"21",X"5E",X"04",X"22",X"54",X"61",
		X"21",X"F7",X"3E",X"AF",X"32",X"52",X"61",X"FB",X"CD",X"18",X"20",X"21",X"38",X"5B",X"22",X"40",
		X"61",X"AF",X"32",X"42",X"61",X"3A",X"52",X"61",X"FE",X"01",X"20",X"F9",X"CD",X"26",X"20",X"DD",
		X"21",X"9C",X"65",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"3E",X"FF",X"DD",X"77",
		X"03",X"AF",X"32",X"58",X"61",X"32",X"C7",X"61",X"3A",X"7D",X"61",X"FE",X"01",X"28",X"14",X"3A",
		X"7C",X"61",X"C6",X"01",X"E6",X"01",X"32",X"7C",X"61",X"3A",X"7D",X"61",X"47",X"FE",X"02",X"78",
		X"CC",X"70",X"2A",X"3A",X"56",X"60",X"FE",X"00",X"20",X"1B",X"3A",X"7C",X"61",X"C6",X"01",X"E6",
		X"01",X"32",X"7C",X"61",X"3A",X"7D",X"61",X"47",X"FE",X"02",X"78",X"CC",X"70",X"2A",X"3A",X"56",
		X"60",X"FE",X"00",X"28",X"67",X"3D",X"32",X"56",X"60",X"CD",X"91",X"35",X"AF",X"32",X"08",X"60",
		X"32",X"4E",X"60",X"32",X"4D",X"60",X"32",X"8F",X"60",X"32",X"77",X"60",X"32",X"37",X"60",X"32",
		X"4F",X"60",X"CD",X"57",X"29",X"3E",X"01",X"C9",X"11",X"BD",X"61",X"01",X"06",X"00",X"ED",X"B0",
		X"3E",X"01",X"32",X"F3",X"61",X"C9",X"DD",X"21",X"44",X"61",X"3E",X"00",X"06",X"06",X"CD",X"54",
		X"20",X"AF",X"32",X"52",X"61",X"32",X"51",X"61",X"32",X"25",X"60",X"32",X"28",X"60",X"32",X"4E",
		X"60",X"32",X"29",X"60",X"32",X"13",X"60",X"32",X"4D",X"60",X"32",X"59",X"61",X"32",X"5E",X"61",
		X"32",X"C7",X"61",X"C9",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F9",X"C9",X"21",X"6E",X"92",X"11",
		X"A1",X"56",X"CD",X"F9",X"30",X"AF",X"32",X"54",X"60",X"06",X"0A",X"21",X"00",X"30",X"2B",X"FB",
		X"3E",X"01",X"32",X"53",X"60",X"32",X"F1",X"61",X"7C",X"FE",X"00",X"20",X"F1",X"10",X"EC",X"CD",
		X"03",X"2D",X"AF",X"32",X"10",X"62",X"3A",X"00",X"60",X"FE",X"00",X"20",X"3C",X"CD",X"03",X"21",
		X"11",X"AC",X"56",X"21",X"5A",X"93",X"CD",X"F9",X"30",X"11",X"E6",X"20",X"21",X"B5",X"93",X"CD",
		X"D9",X"55",X"3E",X"0E",X"21",X"9A",X"98",X"CD",X"05",X"56",X"3E",X"03",X"21",X"55",X"98",X"CD",
		X"05",X"56",X"3E",X"11",X"32",X"B5",X"9B",X"CD",X"8D",X"2F",X"3A",X"B5",X"91",X"FE",X"1F",X"20",
		X"F9",X"3E",X"01",X"32",X"00",X"A0",X"CD",X"34",X"2C",X"F3",X"CD",X"5B",X"35",X"CD",X"67",X"35",
		X"CD",X"63",X"2A",X"AF",X"32",X"53",X"60",X"32",X"F1",X"61",X"3A",X"00",X"60",X"FE",X"00",X"CC",
		X"00",X"37",X"FB",X"3E",X"01",X"C9",X"0E",X"10",X"42",X"59",X"10",X"56",X"41",X"4C",X"41",X"44",
		X"4F",X"4E",X"10",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",X"49",X"4F",X"4E",X"10",X"31",X"39",
		X"38",X"32",X"3F",X"3E",X"00",X"32",X"03",X"A0",X"CD",X"00",X"2A",X"3E",X"30",X"CD",X"EC",X"29",
		X"06",X"01",X"21",X"80",X"65",X"3E",X"00",X"CD",X"F1",X"29",X"CD",X"EC",X"1D",X"3E",X"01",X"32",
		X"03",X"A0",X"C9",X"3A",X"00",X"A0",X"21",X"70",X"59",X"E6",X"03",X"85",X"6F",X"7C",X"CE",X"00",
		X"67",X"7E",X"2A",X"95",X"60",X"77",X"C9",X"3A",X"59",X"61",X"FE",X"01",X"C8",X"3A",X"5E",X"61",
		X"FE",X"01",X"C8",X"0A",X"D9",X"FE",X"00",X"C2",X"A7",X"21",X"2A",X"09",X"60",X"3A",X"0D",X"60",
		X"FD",X"BE",X"02",X"C0",X"FD",X"56",X"01",X"FD",X"5E",X"00",X"D5",X"13",X"13",X"CD",X"45",X"19",
		X"E5",X"AF",X"ED",X"52",X"E1",X"28",X"07",X"CD",X"85",X"35",X"28",X"02",X"D1",X"C9",X"D1",X"CD",
		X"A4",X"19",X"78",X"FE",X"00",X"C8",X"62",X"6B",X"22",X"F6",X"61",X"AF",X"32",X"7E",X"62",X"DD",
		X"21",X"80",X"65",X"FD",X"7E",X"04",X"DD",X"77",X"1C",X"FD",X"7E",X"05",X"DD",X"77",X"1D",X"AF",
		X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",X"7E",X"04",X"FE",X"37",X"20",X"05",X"3E",X"01",X"FD",
		X"77",X"14",X"3E",X"01",X"D9",X"02",X"C9",X"FD",X"7E",X"00",X"FE",X"00",X"C0",X"3A",X"82",X"65",
		X"FE",X"D0",X"D0",X"CD",X"A4",X"19",X"78",X"FE",X"00",X"C8",X"DD",X"21",X"9C",X"65",X"3A",X"0D",
		X"60",X"32",X"98",X"60",X"CD",X"8C",X"55",X"E5",X"3A",X"0D",X"60",X"FD",X"77",X"02",X"CD",X"2D",
		X"22",X"67",X"AF",X"7D",X"D6",X"22",X"6F",X"7C",X"DE",X"00",X"67",X"FD",X"75",X"00",X"FD",X"74",
		X"01",X"3A",X"0D",X"60",X"FD",X"77",X"02",X"C5",X"CD",X"85",X"3C",X"78",X"C1",X"FE",X"00",X"CA",
		X"B7",X"3C",X"E1",X"7E",X"FE",X"E0",X"E5",X"CA",X"B7",X"3C",X"E1",X"E5",X"AF",X"7D",X"D6",X"20",
		X"7C",X"DE",X"00",X"67",X"E1",X"7E",X"FE",X"E0",X"C8",X"D9",X"3A",X"C7",X"61",X"FE",X"01",X"20",
		X"05",X"3E",X"28",X"08",X"18",X"03",X"3E",X"20",X"08",X"AF",X"02",X"FD",X"6E",X"00",X"FD",X"66",
		X"01",X"FD",X"7E",X"06",X"CD",X"17",X"34",X"3E",X"FF",X"32",X"9F",X"65",X"C9",X"FE",X"01",X"20",
		X"04",X"7C",X"C6",X"50",X"C9",X"FE",X"02",X"20",X"04",X"7C",X"C6",X"4C",X"C9",X"7C",X"C6",X"48",
		X"C9",X"FD",X"21",X"56",X"61",X"FD",X"7E",X"00",X"FE",X"01",X"C8",X"3A",X"99",X"60",X"32",X"98",
		X"60",X"DD",X"E5",X"21",X"00",X"05",X"CD",X"90",X"5C",X"21",X"09",X"3F",X"CD",X"18",X"20",X"DD",
		X"E1",X"CD",X"BE",X"3D",X"AF",X"32",X"57",X"60",X"3E",X"21",X"32",X"94",X"65",X"2A",X"38",X"60",
		X"FD",X"21",X"37",X"60",X"DD",X"21",X"94",X"65",X"CD",X"05",X"26",X"C9",X"FD",X"21",X"57",X"61",
		X"FD",X"7E",X"00",X"FE",X"01",X"C8",X"3A",X"9A",X"60",X"32",X"98",X"60",X"DD",X"E5",X"21",X"00",
		X"05",X"CD",X"90",X"5C",X"21",X"09",X"3F",X"CD",X"18",X"20",X"DD",X"E1",X"CD",X"BE",X"3D",X"AF",
		X"32",X"97",X"60",X"3E",X"21",X"32",X"98",X"65",X"2A",X"78",X"60",X"FD",X"21",X"77",X"60",X"DD",
		X"21",X"98",X"65",X"CD",X"05",X"26",X"C9",X"C5",X"FD",X"E5",X"DD",X"E5",X"06",X"03",X"DD",X"21",
		X"CC",X"61",X"DD",X"7E",X"00",X"08",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"08",X"FD",X"77",X"00",
		X"DD",X"23",X"FD",X"23",X"10",X"EC",X"DD",X"E1",X"FD",X"E1",X"C1",X"C9",X"DD",X"21",X"9C",X"60",
		X"3E",X"04",X"32",X"7A",X"62",X"06",X"13",X"DD",X"E5",X"C5",X"CD",X"51",X"31",X"C1",X"DD",X"E1",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"3E",X"01",X"32",X"7A",X"62",X"10",X"EA",X"3A",X"C7",X"61",
		X"FE",X"01",X"28",X"1C",X"3A",X"0D",X"60",X"47",X"FD",X"21",X"C4",X"61",X"FD",X"7E",X"02",X"B8",
		X"20",X"0E",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"3E",X"28",X"08",X"3E",X"EC",X"CD",X"17",X"34",
		X"3A",X"0D",X"60",X"47",X"FD",X"21",X"CC",X"61",X"FD",X"7E",X"02",X"B8",X"20",X"22",X"FD",X"6E",
		X"00",X"FD",X"66",X"01",X"7E",X"CD",X"73",X"35",X"20",X"16",X"E5",X"D5",X"11",X"20",X"00",X"19",
		X"7E",X"CD",X"73",X"35",X"D1",X"E1",X"20",X"08",X"3E",X"20",X"08",X"3E",X"E4",X"CD",X"17",X"34",
		X"06",X"04",X"FD",X"21",X"D3",X"61",X"11",X"CC",X"61",X"C5",X"FD",X"E5",X"D5",X"CD",X"B7",X"22",
		X"1A",X"6F",X"13",X"1A",X"67",X"1B",X"3A",X"0D",X"60",X"FD",X"E1",X"FD",X"BE",X"02",X"FD",X"E5",
		X"20",X"1C",X"7E",X"CD",X"73",X"35",X"20",X"16",X"E5",X"D5",X"11",X"20",X"00",X"19",X"7E",X"CD",
		X"73",X"35",X"D1",X"E1",X"20",X"08",X"3E",X"20",X"08",X"3E",X"E4",X"CD",X"17",X"34",X"D1",X"FD",
		X"E1",X"C1",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"BF",X"C9",X"10",X"BF",X"C9",X"90",X"49",
		X"A0",X"C4",X"20",X"5C",X"02",X"4C",X"05",X"7C",X"00",X"46",X"20",X"48",X"90",X"C0",X"81",X"41",
		X"22",X"49",X"80",X"40",X"00",X"42",X"10",X"48",X"10",X"47",X"10",X"41",X"00",X"5D",X"00",X"46",
		X"11",X"41",X"00",X"D4",X"10",X"44",X"10",X"48",X"33",X"46",X"20",X"CC",X"20",X"4E",X"00",X"6A",
		X"02",X"4A",X"10",X"4D",X"05",X"48",X"20",X"60",X"34",X"42",X"08",X"C0",X"23",X"56",X"A2",X"4D",
		X"10",X"40",X"90",X"4A",X"10",X"4B",X"12",X"4A",X"A0",X"44",X"00",X"DC",X"10",X"C2",X"B8",X"6F",
		X"00",X"48",X"30",X"4E",X"A4",X"44",X"00",X"48",X"22",X"46",X"00",X"47",X"28",X"4D",X"00",X"42",
		X"E7",X"9E",X"06",X"A0",X"C6",X"99",X"C0",X"A3",X"54",X"B4",X"42",X"A3",X"74",X"3E",X"9E",X"12",
		X"5E",X"A8",X"23",X"10",X"42",X"11",X"6F",X"30",X"40",X"3D",X"D3",X"22",X"A2",X"39",X"C1",X"10",
		X"43",X"32",X"61",X"9A",X"41",X"22",X"09",X"10",X"42",X"15",X"83",X"38",X"26",X"BB",X"8D",X"3B",
		X"41",X"3C",X"E2",X"05",X"C2",X"AB",X"C2",X"34",X"CC",X"B0",X"6B",X"12",X"C7",X"AB",X"83",X"0E",
		X"86",X"2E",X"52",X"11",X"E0",X"24",X"08",X"B3",X"8B",X"10",X"8E",X"30",X"DC",X"0D",X"98",X"A2",
		X"EC",X"9A",X"00",X"04",X"CD",X"15",X"CF",X"06",X"4E",X"98",X"86",X"B0",X"4D",X"09",X"C6",X"13",
		X"81",X"92",X"0C",X"B3",X"40",X"92",X"C3",X"95",X"D2",X"11",X"D3",X"18",X"56",X"2D",X"02",X"1E",
		X"37",X"28",X"64",X"81",X"62",X"9A",X"CF",X"B5",X"56",X"BA",X"C1",X"2F",X"D9",X"91",X"87",X"BA",
		X"C3",X"CB",X"29",X"C3",X"DC",X"29",X"31",X"F0",X"67",X"3E",X"3F",X"CD",X"EC",X"29",X"CD",X"00",
		X"2A",X"3E",X"01",X"32",X"03",X"A0",X"21",X"96",X"36",X"11",X"17",X"62",X"01",X"50",X"00",X"ED",
		X"B0",X"C3",X"1C",X"12",X"3A",X"10",X"62",X"FE",X"01",X"20",X"3E",X"3A",X"6D",X"62",X"FE",X"20",
		X"DC",X"BD",X"24",X"FE",X"30",X"DC",X"F2",X"24",X"AF",X"32",X"6D",X"62",X"C9",X"3A",X"6E",X"62",
		X"FE",X"01",X"28",X"13",X"CD",X"01",X"25",X"28",X"10",X"11",X"5A",X"57",X"CD",X"F9",X"30",X"CD",
		X"E9",X"24",X"3E",X"01",X"32",X"6E",X"62",X"F1",X"C9",X"11",X"63",X"57",X"CD",X"F9",X"30",X"CD",
		X"E9",X"24",X"3E",X"01",X"32",X"6E",X"62",X"F1",X"C9",X"3E",X"02",X"21",X"40",X"98",X"CD",X"05",
		X"56",X"C9",X"CD",X"01",X"25",X"11",X"6C",X"57",X"CD",X"F9",X"30",X"AF",X"32",X"6E",X"62",X"F1",
		X"C9",X"3A",X"7C",X"61",X"21",X"A0",X"93",X"FE",X"01",X"C0",X"21",X"20",X"91",X"C9",X"2B",X"CD",
		X"C8",X"25",X"23",X"CD",X"C8",X"25",X"C9",X"3A",X"0D",X"60",X"FE",X"02",X"C0",X"3A",X"83",X"65",
		X"FE",X"C0",X"C0",X"3A",X"82",X"65",X"FE",X"40",X"C0",X"3A",X"CF",X"61",X"FE",X"00",X"C8",X"3A",
		X"9C",X"65",X"FE",X"B8",X"28",X"03",X"FE",X"B7",X"C0",X"3A",X"18",X"93",X"FE",X"E0",X"C8",X"FE",
		X"E6",X"C8",X"FE",X"E4",X"C8",X"FE",X"D0",X"C8",X"3A",X"18",X"93",X"FE",X"02",X"28",X"0B",X"3D",
		X"3D",X"32",X"18",X"93",X"3D",X"32",X"19",X"93",X"18",X"08",X"3E",X"E0",X"32",X"18",X"93",X"32",
		X"19",X"93",X"3A",X"18",X"93",X"32",X"7D",X"62",X"C9",X"C5",X"E5",X"D5",X"AF",X"32",X"0B",X"60",
		X"11",X"FA",X"46",X"ED",X"52",X"20",X"0A",X"CD",X"A1",X"25",X"28",X"05",X"3E",X"02",X"32",X"0B",
		X"60",X"D1",X"E1",X"C1",X"C9",X"C5",X"E5",X"D5",X"AF",X"32",X"0B",X"60",X"11",X"3A",X"47",X"ED",
		X"52",X"20",X"0A",X"CD",X"A1",X"25",X"28",X"05",X"3E",X"02",X"32",X"0B",X"60",X"D1",X"E1",X"C1",
		X"C9",X"21",X"18",X"93",X"7E",X"21",X"AE",X"25",X"01",X"05",X"00",X"ED",X"B1",X"C9",X"0A",X"08",
		X"06",X"04",X"02",X"3A",X"0D",X"60",X"FE",X"02",X"C0",X"3A",X"E8",X"61",X"FE",X"20",X"C0",X"E5",
		X"21",X"0F",X"57",X"7E",X"FE",X"44",X"E1",X"C8",X"7E",X"FD",X"21",X"FC",X"25",X"11",X"EB",X"25",
		X"4F",X"06",X"07",X"1A",X"B9",X"28",X"06",X"13",X"FD",X"23",X"10",X"F7",X"C9",X"DD",X"7E",X"03",
		X"E6",X"F0",X"47",X"FD",X"7E",X"00",X"B0",X"DD",X"77",X"03",X"C9",X"F1",X"F2",X"F3",X"F4",X"F5",
		X"F6",X"F7",X"FB",X"F6",X"FF",X"F7",X"F6",X"F5",X"F4",X"F3",X"F2",X"F1",X"02",X"03",X"04",X"05",
		X"06",X"07",X"08",X"08",X"08",X"CD",X"40",X"26",X"78",X"32",X"0C",X"60",X"FE",X"00",X"C8",X"FD",
		X"7E",X"00",X"FE",X"01",X"C8",X"7E",X"4F",X"11",X"F4",X"25",X"06",X"08",X"1A",X"B9",X"C8",X"13",
		X"10",X"FA",X"3A",X"0C",X"60",X"FE",X"05",X"30",X"09",X"47",X"DD",X"7E",X"03",X"90",X"DD",X"77",
		X"03",X"C9",X"2F",X"E6",X"07",X"C6",X"01",X"47",X"DD",X"7E",X"03",X"80",X"DD",X"77",X"03",X"C9",
		X"DD",X"7E",X"03",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"06",X"00",X"CB",
		X"07",X"CB",X"10",X"CB",X"07",X"CB",X"10",X"CB",X"07",X"CB",X"10",X"CD",X"23",X"29",X"C9",X"CD",
		X"16",X"2A",X"3E",X"3F",X"CD",X"EC",X"29",X"3A",X"00",X"B8",X"21",X"00",X"48",X"11",X"00",X"90",
		X"01",X"00",X"04",X"ED",X"B0",X"21",X"44",X"9B",X"06",X"04",X"CD",X"7B",X"29",X"21",X"24",X"99",
		X"06",X"0F",X"CD",X"7B",X"29",X"21",X"44",X"98",X"06",X"04",X"CD",X"7B",X"29",X"21",X"71",X"98",
		X"06",X"03",X"CD",X"7B",X"29",X"21",X"31",X"99",X"06",X"04",X"CD",X"7B",X"29",X"21",X"50",X"9B",
		X"06",X"04",X"CD",X"7B",X"29",X"21",X"58",X"9B",X"06",X"04",X"CD",X"7B",X"29",X"21",X"18",X"9A",
		X"06",X"08",X"CD",X"7B",X"29",X"21",X"B4",X"99",X"06",X"0B",X"CD",X"7B",X"29",X"21",X"D8",X"98",
		X"06",X"07",X"CD",X"7B",X"29",X"21",X"C8",X"98",X"06",X"0A",X"CD",X"7B",X"29",X"21",X"9B",X"98",
		X"06",X"1A",X"CD",X"85",X"29",X"21",X"25",X"99",X"CD",X"89",X"29",X"21",X"85",X"9A",X"CD",X"89",
		X"29",X"21",X"45",X"9B",X"CD",X"89",X"29",X"21",X"59",X"9B",X"CD",X"89",X"29",X"21",X"19",X"9A",
		X"CD",X"89",X"29",X"21",X"D9",X"9A",X"CD",X"89",X"29",X"21",X"B5",X"9A",X"CD",X"89",X"29",X"21",
		X"51",X"9B",X"CD",X"89",X"29",X"21",X"D9",X"98",X"CD",X"89",X"29",X"21",X"79",X"99",X"CD",X"89",
		X"29",X"21",X"15",X"9A",X"CD",X"89",X"29",X"21",X"29",X"99",X"CD",X"89",X"29",X"21",X"C9",X"99",
		X"CD",X"89",X"29",X"21",X"B8",X"9A",X"3E",X"3F",X"77",X"11",X"05",X"57",X"21",X"40",X"92",X"CD",
		X"F9",X"30",X"21",X"84",X"65",X"3E",X"33",X"77",X"23",X"3E",X"0C",X"77",X"23",X"3E",X"2F",X"77",
		X"23",X"3A",X"00",X"B8",X"3A",X"66",X"61",X"77",X"CD",X"26",X"1E",X"CD",X"10",X"31",X"CD",X"EB",
		X"3D",X"C0",X"21",X"00",X"52",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"C9",X"CD",X"16",X"2A",
		X"3E",X"3F",X"CD",X"EC",X"29",X"3A",X"00",X"B8",X"21",X"00",X"44",X"11",X"00",X"90",X"01",X"00",
		X"04",X"ED",X"B0",X"21",X"B0",X"99",X"06",X"11",X"CD",X"7B",X"29",X"21",X"0B",X"9A",X"06",X"0A",
		X"CD",X"7B",X"29",X"21",X"07",X"9B",X"06",X"06",X"CD",X"7B",X"29",X"21",X"5B",X"99",X"06",X"08",
		X"CD",X"7B",X"29",X"21",X"BB",X"9A",X"06",X"09",X"CD",X"7B",X"29",X"21",X"A7",X"99",X"06",X"08",
		X"CD",X"7B",X"29",X"21",X"44",X"98",X"06",X"08",X"CD",X"7B",X"29",X"21",X"50",X"98",X"06",X"09",
		X"CD",X"7B",X"29",X"21",X"58",X"98",X"06",X"04",X"CD",X"7B",X"29",X"21",X"AA",X"99",X"06",X"0D",
		X"CD",X"85",X"29",X"21",X"5B",X"98",X"06",X"05",X"CD",X"85",X"29",X"21",X"9E",X"98",X"06",X"1A",
		X"CD",X"85",X"29",X"21",X"AA",X"9B",X"3E",X"2F",X"77",X"21",X"31",X"99",X"CD",X"89",X"29",X"21",
		X"C5",X"98",X"CD",X"89",X"29",X"21",X"FC",X"9A",X"CD",X"89",X"29",X"21",X"28",X"9A",X"CD",X"89",
		X"29",X"21",X"D1",X"99",X"CD",X"89",X"29",X"21",X"5C",X"99",X"CD",X"89",X"29",X"21",X"1C",X"9A",
		X"CD",X"89",X"29",X"21",X"EC",X"9A",X"CD",X"89",X"29",X"21",X"08",X"9B",X"CD",X"89",X"29",X"21",
		X"91",X"9B",X"CD",X"89",X"29",X"21",X"FB",X"99",X"3E",X"3F",X"77",X"21",X"07",X"9A",X"77",X"21",
		X"98",X"98",X"77",X"3A",X"00",X"B8",X"11",X"05",X"57",X"21",X"40",X"92",X"CD",X"F9",X"30",X"21",
		X"84",X"65",X"3E",X"33",X"77",X"3E",X"04",X"23",X"77",X"3E",X"97",X"23",X"77",X"3A",X"65",X"61",
		X"23",X"77",X"3A",X"00",X"B8",X"CD",X"26",X"1E",X"CD",X"10",X"31",X"C9",X"CD",X"16",X"2A",X"3E",
		X"3F",X"CD",X"EC",X"29",X"3A",X"00",X"B8",X"21",X"00",X"40",X"11",X"00",X"90",X"01",X"00",X"04",
		X"ED",X"B0",X"21",X"07",X"99",X"06",X"0E",X"CD",X"7B",X"29",X"21",X"17",X"99",X"06",X"0E",X"CD",
		X"7B",X"29",X"21",X"5B",X"98",X"06",X"14",X"CD",X"7B",X"29",X"21",X"47",X"98",X"06",X"03",X"CD",
		X"7B",X"29",X"21",X"50",X"98",X"06",X"03",X"CD",X"7B",X"29",X"21",X"3B",X"9B",X"06",X"03",X"CD",
		X"7B",X"29",X"21",X"4A",X"9B",X"06",X"03",X"CD",X"7B",X"29",X"21",X"4A",X"98",X"06",X"03",X"CD",
		X"85",X"29",X"21",X"0A",X"99",X"06",X"0E",X"CD",X"85",X"29",X"21",X"5E",X"98",X"06",X"1A",X"CD",
		X"85",X"29",X"21",X"68",X"9A",X"CD",X"89",X"29",X"21",X"68",X"99",X"CD",X"89",X"29",X"21",X"18",
		X"99",X"CD",X"89",X"29",X"21",X"98",X"99",X"CD",X"89",X"29",X"21",X"78",X"9A",X"CD",X"89",X"29",
		X"21",X"9C",X"98",X"CD",X"89",X"29",X"21",X"9C",X"9A",X"CD",X"89",X"29",X"21",X"71",X"98",X"CD",
		X"89",X"29",X"21",X"3C",X"9B",X"CD",X"89",X"29",X"3E",X"3F",X"21",X"7B",X"9A",X"77",X"21",X"DB",
		X"98",X"77",X"21",X"27",X"9A",X"77",X"21",X"67",X"98",X"77",X"AF",X"21",X"84",X"65",X"77",X"23",
		X"77",X"23",X"77",X"23",X"77",X"3A",X"00",X"B8",X"CD",X"26",X"1E",X"CD",X"10",X"31",X"3A",X"10",
		X"62",X"FE",X"00",X"C8",X"CD",X"EB",X"3D",X"C0",X"21",X"00",X"50",X"22",X"40",X"61",X"AF",X"32",
		X"42",X"61",X"C9",X"3A",X"0D",X"60",X"FE",X"03",X"C0",X"3A",X"97",X"65",X"FE",X"28",X"C0",X"DD",
		X"E5",X"E5",X"D5",X"DD",X"21",X"0C",X"57",X"DD",X"7E",X"00",X"21",X"94",X"29",X"BE",X"C4",X"46",
		X"29",X"D1",X"E1",X"DD",X"E1",X"C9",X"11",X"A9",X"29",X"21",X"E2",X"92",X"C5",X"F5",X"3E",X"07",
		X"08",X"CD",X"F0",X"55",X"F1",X"C1",X"C9",X"3E",X"01",X"32",X"1A",X"60",X"32",X"1B",X"60",X"3E",
		X"80",X"32",X"27",X"60",X"3E",X"40",X"32",X"67",X"60",X"21",X"95",X"29",X"3A",X"00",X"B8",X"11",
		X"88",X"65",X"01",X"14",X"00",X"ED",X"B0",X"CD",X"E0",X"1E",X"C9",X"3E",X"1F",X"11",X"20",X"00",
		X"77",X"19",X"10",X"FC",X"C9",X"3E",X"2F",X"18",X"F4",X"11",X"20",X"00",X"3E",X"1F",X"77",X"19",
		X"77",X"23",X"77",X"C9",X"41",X"35",X"04",X"5F",X"00",X"35",X"04",X"5F",X"00",X"35",X"04",X"D8",
		X"00",X"20",X"0C",X"D0",X"10",X"20",X"0C",X"D0",X"10",X"26",X"11",X"1C",X"11",X"14",X"1F",X"1E",
		X"10",X"11",X"25",X"24",X"1F",X"1D",X"11",X"24",X"19",X"1F",X"1E",X"3F",X"C5",X"01",X"E0",X"FF",
		X"77",X"09",X"C1",X"10",X"F7",X"C9",X"77",X"23",X"10",X"FC",X"C9",X"06",X"08",X"21",X"00",X"60",
		X"AF",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",X"C3",X"83",X"24",X"06",X"08",X"21",X"00",
		X"60",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",X"C3",X"86",X"24",X"06",X"08",X"21",X"00",
		X"98",X"0E",X"00",X"77",X"23",X"F5",X"3A",X"00",X"B8",X"F1",X"0D",X"20",X"F6",X"10",X"F2",X"C9",
		X"06",X"04",X"3E",X"E0",X"21",X"00",X"90",X"0E",X"00",X"77",X"23",X"F5",X"3A",X"00",X"B8",X"F1",
		X"0D",X"20",X"F6",X"10",X"F2",X"C9",X"3E",X"E0",X"3E",X"E0",X"21",X"E4",X"93",X"06",X"1B",X"E5",
		X"C5",X"06",X"20",X"CD",X"BC",X"29",X"C1",X"E1",X"23",X"10",X"F4",X"C9",X"3E",X"00",X"32",X"03",
		X"A0",X"06",X"04",X"3E",X"E0",X"21",X"00",X"90",X"CD",X"07",X"2A",X"3E",X"3F",X"CD",X"EC",X"29",
		X"3A",X"8C",X"62",X"FE",X"01",X"28",X"09",X"11",X"C3",X"56",X"21",X"AF",X"93",X"CD",X"F9",X"30",
		X"06",X"01",X"21",X"80",X"65",X"3E",X"00",X"CD",X"F1",X"29",X"CD",X"10",X"31",X"3E",X"01",X"32",
		X"03",X"A0",X"C9",X"DD",X"21",X"76",X"61",X"06",X"07",X"AF",X"00",X"DD",X"23",X"10",X"FB",X"C9",
		X"3A",X"63",X"61",X"E6",X"80",X"FE",X"00",X"28",X"0C",X"3A",X"7C",X"61",X"2F",X"E6",X"01",X"32",
		X"01",X"A0",X"32",X"02",X"A0",X"DD",X"21",X"9C",X"60",X"FD",X"21",X"7F",X"61",X"06",X"36",X"CD",
		X"BC",X"2A",X"DD",X"21",X"C4",X"61",X"FD",X"21",X"FA",X"61",X"06",X"03",X"CD",X"BC",X"2A",X"3A",
		X"56",X"60",X"F5",X"3A",X"7E",X"61",X"32",X"56",X"60",X"F1",X"32",X"7E",X"61",X"3A",X"90",X"62",
		X"F5",X"3A",X"7D",X"62",X"32",X"90",X"62",X"F1",X"32",X"7D",X"62",X"C9",X"DD",X"7E",X"00",X"F5",
		X"FD",X"7E",X"00",X"DD",X"77",X"00",X"F1",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"10",X"EC",
		X"C9",X"0E",X"0B",X"06",X"07",X"DD",X"7E",X"03",X"C6",X"03",X"91",X"FD",X"BE",X"03",X"28",X"06",
		X"0C",X"10",X"F2",X"3E",X"00",X"C9",X"DD",X"7E",X"02",X"C6",X"08",X"FD",X"BE",X"02",X"38",X"F3",
		X"D6",X"0F",X"FD",X"BE",X"02",X"30",X"EC",X"3E",X"01",X"C9",X"3A",X"98",X"60",X"47",X"3A",X"0D",
		X"60",X"B8",X"C2",X"1E",X"2C",X"E5",X"FD",X"E5",X"FD",X"21",X"D3",X"2C",X"FD",X"7E",X"00",X"67",
		X"FD",X"7E",X"01",X"6F",X"AF",X"ED",X"52",X"28",X"18",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",
		X"7E",X"02",X"FE",X"FF",X"20",X"E6",X"2A",X"46",X"61",X"AF",X"77",X"FD",X"E1",X"E1",X"C3",X"84",
		X"2B",X"3E",X"01",X"2A",X"46",X"61",X"7E",X"FE",X"00",X"C2",X"2B",X"2B",X"CD",X"D1",X"2B",X"FD",
		X"E1",X"47",X"FD",X"7E",X"03",X"B8",X"CA",X"C6",X"2B",X"2A",X"46",X"61",X"23",X"23",X"23",X"23",
		X"3E",X"01",X"77",X"E1",X"D5",X"11",X"1C",X"00",X"19",X"D1",X"AF",X"77",X"DD",X"7E",X"07",X"3D",
		X"FD",X"BE",X"03",X"28",X"0C",X"3D",X"FD",X"BE",X"03",X"28",X"06",X"2A",X"95",X"60",X"AF",X"77",
		X"C9",X"DD",X"7E",X"06",X"2A",X"95",X"60",X"FD",X"BE",X"02",X"30",X"04",X"3E",X"40",X"77",X"C9",
		X"3E",X"80",X"77",X"C9",X"7E",X"FE",X"01",X"28",X"09",X"2A",X"46",X"61",X"23",X"23",X"23",X"23",
		X"77",X"C9",X"2A",X"46",X"61",X"3E",X"01",X"77",X"CD",X"D1",X"2B",X"47",X"FD",X"7E",X"03",X"B8",
		X"28",X"25",X"23",X"23",X"23",X"23",X"3E",X"01",X"77",X"3A",X"98",X"60",X"FE",X"02",X"20",X"07",
		X"3E",X"98",X"FD",X"77",X"02",X"18",X"09",X"FE",X"03",X"20",X"05",X"3E",X"30",X"FD",X"77",X"02",
		X"2A",X"95",X"60",X"AF",X"77",X"C9",X"E1",X"2A",X"46",X"61",X"23",X"23",X"23",X"23",X"AF",X"77",
		X"C9",X"3A",X"98",X"60",X"FE",X"03",X"28",X"16",X"FE",X"02",X"C0",X"DD",X"7E",X"03",X"FE",X"80",
		X"3E",X"88",X"D0",X"DD",X"7E",X"02",X"FE",X"98",X"3E",X"40",X"D8",X"3E",X"69",X"C9",X"DD",X"7E",
		X"02",X"FE",X"28",X"06",X"40",X"38",X"02",X"06",X"80",X"DD",X"7E",X"03",X"FE",X"78",X"3E",X"29",
		X"38",X"15",X"DD",X"7E",X"03",X"FE",X"A0",X"3E",X"71",X"38",X"0C",X"DD",X"7E",X"03",X"FE",X"C0",
		X"3E",X"A9",X"38",X"03",X"3E",X"C8",X"C9",X"E5",X"2A",X"95",X"60",X"70",X"E1",X"C9",X"2A",X"46",
		X"61",X"23",X"23",X"23",X"23",X"AF",X"77",X"C9",X"3A",X"78",X"61",X"FE",X"06",X"C0",X"3A",X"A3",
		X"58",X"FE",X"4C",X"C8",X"21",X"00",X"05",X"FB",X"06",X"FF",X"3A",X"00",X"60",X"FE",X"00",X"C0",
		X"3A",X"00",X"B8",X"FB",X"10",X"F4",X"2B",X"7C",X"FE",X"00",X"C8",X"18",X"EB",X"3A",X"ED",X"61",
		X"FE",X"01",X"3E",X"00",X"28",X"22",X"3A",X"78",X"61",X"47",X"3A",X"7C",X"61",X"FE",X"01",X"20",
		X"04",X"3A",X"7B",X"61",X"47",X"3A",X"00",X"B0",X"CB",X"1F",X"CB",X"1F",X"CB",X"1F",X"2F",X"E6",
		X"03",X"80",X"06",X"00",X"CD",X"7C",X"2C",X"78",X"32",X"64",X"61",X"C9",X"FE",X"01",X"D8",X"06",
		X"02",X"FE",X"02",X"D8",X"06",X"04",X"FE",X"03",X"D8",X"06",X"05",X"FE",X"04",X"D8",X"06",X"09",
		X"FE",X"05",X"D8",X"06",X"0A",X"C9",X"DD",X"21",X"94",X"65",X"FD",X"21",X"9C",X"65",X"CD",X"D1",
		X"2A",X"FE",X"01",X"20",X"0F",X"3A",X"58",X"61",X"FE",X"01",X"28",X"08",X"3E",X"01",X"32",X"37",
		X"60",X"32",X"08",X"62",X"DD",X"21",X"98",X"65",X"FD",X"21",X"9C",X"65",X"CD",X"D1",X"2A",X"FE",
		X"01",X"20",X"0F",X"3A",X"58",X"61",X"FE",X"01",X"28",X"08",X"3E",X"01",X"32",X"77",X"60",X"32",
		X"09",X"62",X"C9",X"45",X"44",X"40",X"45",X"4F",X"40",X"45",X"53",X"40",X"45",X"A4",X"80",X"45",
		X"AA",X"80",X"45",X"B3",X"80",X"4A",X"E4",X"40",X"4A",X"E7",X"40",X"4A",X"F0",X"40",X"4A",X"F7",
		X"40",X"4A",X"FB",X"40",X"4B",X"44",X"80",X"4B",X"47",X"80",X"4B",X"53",X"80",X"4B",X"5B",X"80",
		X"FF",X"FF",X"FF",X"3A",X"10",X"62",X"FE",X"01",X"C0",X"FD",X"21",X"76",X"61",X"CD",X"D8",X"2D",
		X"78",X"FE",X"05",X"38",X"0B",X"FD",X"21",X"79",X"61",X"CD",X"D8",X"2D",X"78",X"FE",X"05",X"D0",
		X"CD",X"03",X"21",X"CD",X"FB",X"2F",X"3A",X"6C",X"62",X"FE",X"01",X"CC",X"70",X"2A",X"CD",X"8D",
		X"2F",X"3E",X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",X"FD",X"21",X"76",X"61",X"CD",X"D8",X"2D",
		X"78",X"FE",X"05",X"D2",X"71",X"2D",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"D5",X"11",X"F0",X"FF",
		X"DD",X"19",X"D1",X"DD",X"E5",X"23",X"23",X"E5",X"CD",X"04",X"2E",X"3E",X"60",X"32",X"E8",X"61",
		X"E1",X"CD",X"8D",X"2F",X"DD",X"E1",X"3E",X"01",X"32",X"79",X"62",X"CD",X"58",X"2E",X"CD",X"8D",
		X"2F",X"3A",X"7D",X"61",X"FE",X"01",X"28",X"5B",X"3A",X"00",X"B0",X"E6",X"80",X"FE",X"80",X"28",
		X"08",X"3E",X"00",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3A",X"26",X"60",X"E6",X"80",X"FE",X"80",
		X"28",X"F7",X"FD",X"21",X"79",X"61",X"CD",X"D8",X"2D",X"78",X"FE",X"05",X"30",X"35",X"CD",X"8D",
		X"2F",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"D5",X"11",X"F0",X"FF",X"DD",X"19",X"D1",X"DD",X"E5",
		X"23",X"23",X"E5",X"CD",X"04",X"2E",X"3E",X"60",X"32",X"E8",X"61",X"E1",X"CD",X"8D",X"2F",X"DD",
		X"E1",X"3E",X"00",X"32",X"79",X"62",X"CD",X"19",X"2F",X"CD",X"19",X"2F",X"CD",X"19",X"2F",X"CD",
		X"58",X"2E",X"C9",X"AF",X"32",X"67",X"62",X"C9",X"DD",X"21",X"17",X"62",X"11",X"10",X"00",X"21",
		X"0F",X"92",X"06",X"05",X"FD",X"7E",X"02",X"DD",X"BE",X"02",X"D8",X"20",X"10",X"FD",X"7E",X"01",
		X"DD",X"BE",X"01",X"D8",X"20",X"07",X"FD",X"7E",X"00",X"DD",X"BE",X"00",X"D8",X"DD",X"19",X"2B",
		X"2B",X"10",X"E1",X"C9",X"C5",X"DD",X"21",X"17",X"62",X"78",X"FE",X"04",X"30",X"11",X"C5",X"06",
		X"10",X"DD",X"7E",X"10",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F6",X"C1",X"04",X"18",X"EA",X"C1",
		X"DD",X"21",X"17",X"62",X"78",X"FE",X"04",X"30",X"05",X"DD",X"19",X"04",X"18",X"F6",X"FD",X"7E",
		X"00",X"DD",X"77",X"00",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"FD",X"7E",X"02",X"DD",X"77",X"02",
		X"C5",X"06",X"0D",X"DD",X"E5",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"3E",X"10",X"DD",X"77",X"00",
		X"DD",X"23",X"10",X"F9",X"DD",X"E1",X"C1",X"C9",X"06",X"11",X"3E",X"00",X"32",X"78",X"62",X"3A",
		X"79",X"62",X"FE",X"01",X"20",X"05",X"CD",X"9C",X"30",X"18",X"0C",X"3A",X"00",X"B0",X"E6",X"80",
		X"FE",X"80",X"28",X"F2",X"CD",X"B8",X"30",X"3A",X"78",X"62",X"E6",X"10",X"FE",X"10",X"CC",X"B2",
		X"2E",X"3A",X"78",X"62",X"E6",X"08",X"FE",X"08",X"CC",X"C1",X"2E",X"3A",X"78",X"62",X"E6",X"40",
		X"FE",X"40",X"CC",X"D0",X"2E",X"3A",X"78",X"62",X"E6",X"20",X"FE",X"20",X"CC",X"EE",X"2E",X"3A",
		X"78",X"62",X"E6",X"80",X"FE",X"80",X"C8",X"3A",X"E8",X"61",X"FE",X"00",X"C8",X"CD",X"0A",X"2F",
		X"18",X"AD",X"78",X"FE",X"29",X"20",X"02",X"06",X"10",X"04",X"CD",X"0A",X"2F",X"CD",X"19",X"2F",
		X"C9",X"78",X"FE",X"10",X"20",X"02",X"06",X"2A",X"05",X"CD",X"0A",X"2F",X"CD",X"19",X"2F",X"C9",
		X"7D",X"E6",X"F0",X"FE",X"00",X"20",X"04",X"7C",X"FE",X"92",X"C8",X"06",X"10",X"CD",X"0A",X"2F",
		X"11",X"20",X"00",X"19",X"DD",X"2B",X"46",X"CD",X"0A",X"2F",X"CD",X"19",X"2F",X"C9",X"7D",X"E6",
		X"F0",X"FE",X"80",X"20",X"04",X"7C",X"FE",X"90",X"C8",X"11",X"20",X"00",X"AF",X"ED",X"52",X"DD",
		X"23",X"06",X"11",X"CD",X"0A",X"2F",X"CD",X"19",X"2F",X"C9",X"78",X"DD",X"77",X"00",X"77",X"E5",
		X"7C",X"C6",X"08",X"67",X"3E",X"04",X"77",X"E1",X"C9",X"C5",X"F5",X"E5",X"06",X"70",X"21",X"00",
		X"03",X"2B",X"7C",X"FE",X"00",X"20",X"FA",X"10",X"F5",X"E1",X"F1",X"C1",X"C9",X"21",X"25",X"93",
		X"11",X"4F",X"57",X"CD",X"F9",X"30",X"21",X"05",X"92",X"11",X"55",X"57",X"CD",X"F9",X"30",X"21",
		X"E3",X"92",X"11",X"90",X"56",X"CD",X"F9",X"30",X"21",X"83",X"98",X"3E",X"0E",X"CD",X"05",X"56",
		X"11",X"00",X"4D",X"21",X"82",X"93",X"3E",X"12",X"08",X"CD",X"F0",X"55",X"11",X"1B",X"4D",X"21",
		X"90",X"93",X"3E",X"12",X"08",X"CD",X"F0",X"55",X"06",X"0D",X"3E",X"8B",X"21",X"83",X"93",X"CD",
		X"7D",X"2F",X"3E",X"8E",X"06",X"0D",X"21",X"63",X"90",X"CD",X"7D",X"2F",X"C9",X"77",X"E5",X"F5",
		X"7C",X"C6",X"08",X"67",X"3E",X"10",X"77",X"F1",X"E1",X"23",X"10",X"F1",X"C9",X"DD",X"E5",X"C5",
		X"E5",X"D5",X"CD",X"2D",X"2F",X"11",X"20",X"00",X"21",X"8F",X"92",X"DD",X"21",X"17",X"62",X"06",
		X"05",X"C5",X"E5",X"06",X"03",X"DD",X"7E",X"00",X"E6",X"0F",X"CD",X"0E",X"2F",X"DD",X"7E",X"00",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"11",X"20",X"00",X"19",X"CD",X"0E",X"2F",X"DD",X"23",X"19",
		X"10",X"E3",X"E1",X"2B",X"2B",X"C1",X"11",X"0D",X"00",X"DD",X"19",X"10",X"D4",X"11",X"20",X"00",
		X"DD",X"21",X"17",X"62",X"21",X"0F",X"92",X"06",X"05",X"C5",X"E5",X"DD",X"23",X"DD",X"23",X"DD",
		X"23",X"06",X"0D",X"DD",X"7E",X"00",X"CD",X"0E",X"2F",X"DD",X"23",X"ED",X"52",X"10",X"F4",X"E1",
		X"2B",X"2B",X"C1",X"10",X"E4",X"D1",X"E1",X"C1",X"DD",X"E1",X"C9",X"3E",X"01",X"32",X"67",X"62",
		X"21",X"72",X"93",X"11",X"1E",X"57",X"CD",X"F9",X"30",X"21",X"73",X"93",X"11",X"37",X"57",X"CD",
		X"F9",X"30",X"21",X"7D",X"93",X"11",X"75",X"57",X"CD",X"F9",X"30",X"11",X"00",X"4D",X"21",X"91",
		X"93",X"3E",X"12",X"08",X"CD",X"F0",X"55",X"11",X"1B",X"4D",X"21",X"9E",X"93",X"3E",X"12",X"08",
		X"CD",X"F0",X"55",X"06",X"0C",X"21",X"92",X"93",X"3E",X"8B",X"CD",X"7D",X"2F",X"06",X"0C",X"3E",
		X"8E",X"21",X"72",X"90",X"CD",X"7D",X"2F",X"11",X"36",X"4D",X"21",X"75",X"92",X"CD",X"DB",X"30",
		X"11",X"4A",X"4D",X"21",X"B8",X"91",X"CD",X"DB",X"30",X"11",X"5E",X"4D",X"21",X"9B",X"92",X"CD",
		X"DB",X"30",X"11",X"72",X"4D",X"21",X"F8",X"92",X"CD",X"DB",X"30",X"11",X"86",X"4D",X"21",X"58",
		X"92",X"CD",X"D4",X"30",X"11",X"8C",X"4D",X"21",X"16",X"92",X"CD",X"D4",X"30",X"11",X"8E",X"4D",
		X"21",X"17",X"92",X"CD",X"D4",X"30",X"11",X"90",X"4D",X"21",X"19",X"92",X"CD",X"D4",X"30",X"11",
		X"92",X"4D",X"21",X"1A",X"92",X"CD",X"D4",X"30",X"CD",X"2D",X"2F",X"C9",X"AF",X"32",X"07",X"A0",
		X"3E",X"07",X"D3",X"08",X"3E",X"38",X"D3",X"09",X"3E",X"0E",X"D3",X"08",X"DB",X"0C",X"2F",X"32",
		X"78",X"62",X"3E",X"01",X"32",X"07",X"A0",X"C9",X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",
		X"3E",X"38",X"D3",X"09",X"3E",X"0F",X"D3",X"08",X"DB",X"0C",X"2F",X"32",X"78",X"62",X"3E",X"01",
		X"32",X"07",X"A0",X"C9",X"3E",X"14",X"08",X"CD",X"F0",X"55",X"C9",X"3E",X"18",X"08",X"CD",X"E5",
		X"30",X"CD",X"F0",X"55",X"C9",X"F5",X"3A",X"00",X"B0",X"E6",X"20",X"FE",X"20",X"20",X"08",X"E5",
		X"EB",X"11",X"0A",X"00",X"19",X"EB",X"E1",X"F1",X"C9",X"F5",X"3A",X"00",X"B0",X"E6",X"20",X"FE",
		X"20",X"28",X"08",X"E5",X"EB",X"11",X"96",X"01",X"19",X"EB",X"E1",X"F1",X"CD",X"D9",X"55",X"C9",
		X"11",X"5A",X"57",X"21",X"A0",X"93",X"CD",X"F9",X"30",X"11",X"63",X"57",X"21",X"20",X"91",X"CD",
		X"F9",X"30",X"C9",X"3A",X"26",X"60",X"FE",X"A5",X"C0",X"11",X"62",X"36",X"21",X"A2",X"93",X"CD",
		X"F0",X"55",X"11",X"7F",X"36",X"21",X"A3",X"93",X"CD",X"F0",X"55",X"18",X"E6",X"DD",X"21",X"CC",
		X"61",X"AF",X"DD",X"77",X"03",X"32",X"E0",X"61",X"32",X"E1",X"61",X"3E",X"FF",X"32",X"9F",X"65",
		X"C9",X"DD",X"7E",X"00",X"6F",X"DD",X"7E",X"01",X"67",X"3A",X"0D",X"60",X"47",X"DD",X"7E",X"02",
		X"B8",X"C0",X"3E",X"D0",X"77",X"E5",X"CD",X"97",X"31",X"E1",X"23",X"7E",X"FE",X"ED",X"28",X"0C",
		X"FE",X"EF",X"28",X"08",X"3E",X"D1",X"77",X"E5",X"CD",X"97",X"31",X"E1",X"11",X"20",X"00",X"19",
		X"7E",X"FE",X"D1",X"C8",X"FE",X"67",X"C8",X"FE",X"27",X"C8",X"FE",X"ED",X"C8",X"FE",X"EF",X"C8",
		X"3E",X"D3",X"77",X"CD",X"97",X"31",X"C9",X"7C",X"FE",X"00",X"C8",X"C6",X"08",X"67",X"3A",X"7A",
		X"62",X"77",X"C9",X"DD",X"21",X"94",X"65",X"3A",X"3B",X"60",X"FE",X"01",X"C8",X"3A",X"56",X"61",
		X"FE",X"01",X"C8",X"3A",X"11",X"62",X"FE",X"01",X"C8",X"CD",X"DF",X"31",X"78",X"32",X"99",X"60",
		X"C9",X"DD",X"21",X"98",X"65",X"3A",X"7B",X"60",X"FE",X"01",X"C8",X"3A",X"57",X"61",X"FE",X"01",
		X"C8",X"3A",X"12",X"62",X"FE",X"01",X"C8",X"CD",X"DF",X"31",X"78",X"32",X"9A",X"60",X"C9",X"3E",
		X"80",X"DD",X"77",X"02",X"3E",X"10",X"DD",X"77",X"03",X"06",X"03",X"3A",X"0D",X"60",X"FE",X"03",
		X"C0",X"06",X"02",X"C9",X"3A",X"F3",X"61",X"FE",X"00",X"C8",X"3C",X"C5",X"47",X"3A",X"75",X"62",
		X"FE",X"01",X"78",X"C1",X"20",X"06",X"FE",X"30",X"20",X"0B",X"18",X"02",X"FE",X"17",X"20",X"05",
		X"3E",X"00",X"32",X"75",X"62",X"32",X"F3",X"61",X"C9",X"3A",X"82",X"65",X"FE",X"E8",X"3E",X"00",
		X"32",X"85",X"62",X"D4",X"43",X"32",X"3A",X"82",X"65",X"FE",X"10",X"DC",X"84",X"32",X"3E",X"00",
		X"32",X"6F",X"62",X"CD",X"FF",X"10",X"F3",X"AF",X"32",X"00",X"A0",X"FB",X"3E",X"01",X"32",X"00",
		X"A0",X"00",X"C9",X"CD",X"74",X"33",X"3A",X"0D",X"60",X"FE",X"01",X"20",X"14",X"CD",X"5D",X"27",
		X"3E",X"11",X"32",X"82",X"65",X"CD",X"E3",X"33",X"CD",X"DC",X"22",X"CD",X"B1",X"33",X"C3",X"CE",
		X"32",X"3A",X"0D",X"60",X"FE",X"02",X"20",X"19",X"3A",X"87",X"65",X"32",X"65",X"61",X"CD",X"5F",
		X"26",X"3E",X"03",X"32",X"0D",X"60",X"CD",X"DC",X"22",X"3E",X"11",X"32",X"82",X"65",X"CD",X"B1",
		X"33",X"C3",X"CE",X"32",X"3E",X"01",X"32",X"85",X"62",X"CD",X"74",X"33",X"3A",X"0D",X"60",X"FE",
		X"01",X"C8",X"FE",X"02",X"20",X"16",X"CD",X"4C",X"28",X"3E",X"01",X"32",X"0D",X"60",X"CD",X"DC",
		X"22",X"3E",X"E3",X"32",X"82",X"65",X"CD",X"B1",X"33",X"C3",X"CE",X"32",X"FE",X"03",X"C0",X"3A",
		X"87",X"65",X"32",X"66",X"61",X"DD",X"21",X"42",X"44",X"DD",X"22",X"81",X"62",X"CD",X"5D",X"27",
		X"3E",X"E3",X"32",X"82",X"65",X"CD",X"E3",X"33",X"CD",X"DC",X"22",X"CD",X"B1",X"33",X"3E",X"01",
		X"32",X"03",X"A0",X"DD",X"21",X"94",X"65",X"FD",X"21",X"80",X"65",X"FD",X"7E",X"03",X"DD",X"BE",
		X"03",X"C2",X"FA",X"32",X"DD",X"7E",X"02",X"FE",X"CD",X"38",X"05",X"CD",X"4E",X"36",X"18",X"0A",
		X"DD",X"7E",X"02",X"FE",X"26",X"30",X"03",X"CD",X"4E",X"36",X"DD",X"21",X"98",X"65",X"FD",X"21",
		X"80",X"65",X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"C2",X"21",X"33",X"DD",X"7E",X"02",X"FE",X"E0",
		X"38",X"05",X"CD",X"58",X"36",X"18",X"0A",X"DD",X"7E",X"02",X"FE",X"10",X"30",X"03",X"CD",X"58",
		X"36",X"3A",X"1C",X"60",X"FE",X"01",X"C8",X"3A",X"1D",X"60",X"FE",X"01",X"C8",X"3A",X"1E",X"60",
		X"FE",X"01",X"C8",X"21",X"83",X"65",X"DD",X"21",X"8C",X"65",X"7E",X"FE",X"40",X"20",X"05",X"CD",
		X"69",X"33",X"18",X"17",X"DD",X"21",X"88",X"65",X"FE",X"E0",X"20",X"05",X"CD",X"69",X"33",X"18",
		X"0A",X"DD",X"21",X"90",X"65",X"FE",X"C8",X"C0",X"CD",X"69",X"33",X"06",X"30",X"C5",X"CD",X"F4",
		X"08",X"C1",X"10",X"F9",X"AF",X"32",X"25",X"60",X"C9",X"DD",X"7E",X"02",X"FE",X"D8",X"D0",X"FE",
		X"18",X"D8",X"F1",X"C9",X"AF",X"32",X"03",X"A0",X"3A",X"C7",X"61",X"FE",X"00",X"CC",X"25",X"1F",
		X"3A",X"59",X"61",X"FE",X"00",X"28",X"0C",X"3A",X"9F",X"65",X"3C",X"32",X"9F",X"65",X"CD",X"83",
		X"16",X"18",X"E1",X"3A",X"3B",X"60",X"FE",X"01",X"20",X"08",X"3E",X"01",X"32",X"EB",X"61",X"32",
		X"3A",X"60",X"3A",X"7B",X"60",X"FE",X"01",X"C0",X"3E",X"01",X"32",X"EC",X"61",X"32",X"7A",X"60",
		X"C9",X"DD",X"21",X"19",X"60",X"21",X"82",X"65",X"FD",X"21",X"8A",X"65",X"11",X"04",X"00",X"CD",
		X"D1",X"33",X"DD",X"23",X"FD",X"19",X"CD",X"D1",X"33",X"DD",X"23",X"FD",X"19",X"CD",X"D1",X"33",
		X"C9",X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"7E",X"FD",X"77",X"00",X"3A",X"0D",X"60",X"3D",X"DD",
		X"77",X"00",X"C9",X"3A",X"7D",X"62",X"32",X"18",X"93",X"FE",X"E0",X"28",X"01",X"3D",X"32",X"19",
		X"93",X"3E",X"02",X"32",X"0D",X"60",X"3E",X"53",X"E5",X"D5",X"C5",X"21",X"B6",X"93",X"11",X"E0",
		X"FF",X"06",X"06",X"77",X"3D",X"F5",X"E5",X"7C",X"C6",X"08",X"67",X"3E",X"1F",X"77",X"E1",X"F1",
		X"19",X"10",X"F0",X"C1",X"D1",X"E1",X"C9",X"C5",X"47",X"7C",X"FE",X"00",X"78",X"C1",X"C8",X"F5",
		X"7E",X"FE",X"D0",X"28",X"06",X"F1",X"CD",X"41",X"34",X"18",X"01",X"F1",X"23",X"3C",X"CD",X"41",
		X"34",X"D5",X"11",X"1F",X"00",X"19",X"D1",X"3C",X"CD",X"41",X"34",X"23",X"3C",X"CD",X"41",X"34",
		X"C9",X"77",X"E5",X"F5",X"7C",X"C6",X"08",X"67",X"08",X"77",X"08",X"F1",X"E1",X"C9",X"3A",X"5E",
		X"61",X"FE",X"01",X"C0",X"DD",X"21",X"94",X"65",X"CD",X"6D",X"34",X"FE",X"01",X"CC",X"41",X"22",
		X"DD",X"21",X"98",X"65",X"CD",X"6D",X"34",X"FE",X"01",X"CC",X"7C",X"22",X"C9",X"FD",X"21",X"9C",
		X"65",X"FD",X"7E",X"02",X"DD",X"BE",X"02",X"28",X"06",X"3C",X"DD",X"BE",X"02",X"20",X"1F",X"FD",
		X"7E",X"03",X"3C",X"3C",X"DD",X"BE",X"03",X"28",X"18",X"3D",X"DD",X"BE",X"03",X"28",X"12",X"3D",
		X"DD",X"BE",X"03",X"28",X"0C",X"3D",X"DD",X"BE",X"03",X"28",X"06",X"3D",X"28",X"03",X"3E",X"00",
		X"C9",X"3E",X"01",X"C9",X"21",X"04",X"A0",X"FD",X"21",X"E5",X"61",X"FD",X"7E",X"00",X"FE",X"00",
		X"28",X"16",X"FD",X"34",X"01",X"FD",X"7E",X"01",X"FE",X"10",X"38",X"0C",X"FE",X"20",X"38",X"0B",
		X"FD",X"35",X"00",X"AF",X"FD",X"77",X"01",X"C9",X"AF",X"77",X"C9",X"3E",X"01",X"77",X"C9",X"3A",
		X"00",X"A0",X"E6",X"3F",X"47",X"00",X"10",X"FD",X"3A",X"00",X"B0",X"E6",X"40",X"FE",X"40",X"3E",
		X"03",X"28",X"02",X"3E",X"04",X"47",X"3A",X"7C",X"61",X"FE",X"01",X"3A",X"78",X"61",X"20",X"03",
		X"3A",X"7B",X"61",X"B8",X"30",X"05",X"AF",X"32",X"86",X"62",X"C9",X"3A",X"86",X"62",X"FE",X"00",
		X"C0",X"3A",X"56",X"60",X"3C",X"32",X"56",X"60",X"3E",X"01",X"32",X"86",X"62",X"C9",X"7E",X"FE",
		X"E0",X"20",X"23",X"3A",X"0D",X"60",X"B8",X"28",X"1D",X"78",X"FE",X"02",X"01",X"65",X"61",X"28",
		X"05",X"FE",X"03",X"01",X"66",X"61",X"0A",X"FE",X"10",X"D8",X"08",X"FE",X"00",X"20",X"03",X"0A",
		X"3D",X"02",X"1A",X"3D",X"12",X"C9",X"AF",X"DD",X"77",X"00",X"FD",X"77",X"00",X"C9",X"21",X"E7",
		X"61",X"7E",X"D6",X"01",X"27",X"77",X"F5",X"23",X"F1",X"7E",X"DE",X"00",X"27",X"77",X"C9",X"11",
		X"9C",X"60",X"21",X"54",X"5C",X"01",X"3A",X"00",X"ED",X"B0",X"C9",X"11",X"9C",X"60",X"21",X"E8",
		X"5A",X"01",X"3A",X"00",X"ED",X"B0",X"C9",X"11",X"7F",X"61",X"21",X"E8",X"5A",X"01",X"3A",X"00",
		X"ED",X"B0",X"C9",X"FE",X"E0",X"C8",X"FE",X"4B",X"C8",X"FE",X"4A",X"C8",X"FE",X"49",X"C8",X"FE",
		X"E4",X"C8",X"FE",X"E6",X"C9",X"E5",X"C5",X"01",X"E0",X"FF",X"09",X"AF",X"ED",X"52",X"C1",X"E1",
		X"C9",X"3A",X"7D",X"61",X"FE",X"01",X"C8",X"3E",X"01",X"32",X"53",X"60",X"32",X"8C",X"62",X"CD",
		X"2C",X"2A",X"11",X"5A",X"57",X"21",X"74",X"92",X"CD",X"F9",X"30",X"11",X"89",X"56",X"21",X"9F",
		X"91",X"CD",X"F9",X"30",X"3A",X"7C",X"61",X"3C",X"32",X"94",X"91",X"3E",X"08",X"21",X"7F",X"98",
		X"CD",X"05",X"56",X"3E",X"00",X"32",X"5F",X"98",X"3E",X"05",X"21",X"41",X"98",X"CD",X"05",X"56",
		X"3E",X"02",X"21",X"40",X"98",X"CD",X"05",X"56",X"21",X"93",X"92",X"11",X"38",X"36",X"3E",X"1F",
		X"08",X"CD",X"F0",X"55",X"21",X"95",X"92",X"11",X"43",X"36",X"3E",X"1F",X"08",X"CD",X"F0",X"55",
		X"3E",X"8E",X"32",X"74",X"91",X"3E",X"8B",X"32",X"94",X"92",X"3E",X"1F",X"32",X"74",X"99",X"32",
		X"94",X"9A",X"CD",X"BE",X"39",X"3E",X"00",X"32",X"03",X"98",X"32",X"07",X"98",X"32",X"0B",X"98",
		X"32",X"0F",X"98",X"32",X"13",X"98",X"32",X"17",X"98",X"32",X"1B",X"98",X"32",X"1F",X"98",X"06",
		X"06",X"21",X"00",X"00",X"2B",X"3A",X"00",X"B8",X"7C",X"FE",X"00",X"20",X"F7",X"10",X"F2",X"3E",
		X"00",X"32",X"53",X"60",X"32",X"8C",X"62",X"C9",X"8A",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"8F",X"3F",X"8C",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8D",X"3F",X"06",X"60",
		X"C5",X"CD",X"6F",X"11",X"C1",X"10",X"F9",X"C9",X"06",X"60",X"C5",X"CD",X"9B",X"11",X"C1",X"10",
		X"F9",X"C9",X"13",X"15",X"10",X"1A",X"15",X"25",X"10",X"1C",X"15",X"10",X"12",X"11",X"17",X"1E",
		X"11",X"22",X"14",X"10",X"11",X"10",X"15",X"24",X"15",X"10",X"13",X"22",X"15",X"15",X"3F",X"20",
		X"11",X"22",X"10",X"26",X"11",X"1C",X"11",X"14",X"1F",X"1E",X"10",X"11",X"25",X"24",X"1F",X"1D",
		X"11",X"24",X"19",X"1F",X"1E",X"3F",X"00",X"42",X"01",X"1A",X"10",X"12",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"51",X"01",X"1A",X"1F",X"1A",X"1F",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"60",X"01",X"20",X"19",X"15",X"22",X"22",X"1F",X"24",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"79",X"01",X"17",X"11",X"23",X"24",X"1F",X"25",X"1E",
		X"15",X"24",X"10",X"10",X"10",X"10",X"00",X"89",X"01",X"16",X"11",X"1E",X"13",X"18",X"1F",X"19",
		X"23",X"10",X"10",X"10",X"10",X"10",X"ED",X"BC",X"FF",X"B5",X"FF",X"85",X"EF",X"B7",X"DF",X"BE",
		X"EF",X"3A",X"7F",X"3F",X"FF",X"25",X"7F",X"B3",X"FF",X"35",X"FF",X"81",X"FF",X"36",X"FF",X"B7",
		X"3E",X"00",X"32",X"03",X"A0",X"CD",X"00",X"2A",X"3E",X"3F",X"CD",X"EC",X"29",X"CD",X"EC",X"1D",
		X"3E",X"01",X"32",X"0D",X"60",X"32",X"03",X"A0",X"32",X"98",X"60",X"32",X"99",X"60",X"32",X"9A",
		X"60",X"AF",X"32",X"08",X"60",X"32",X"37",X"60",X"32",X"4E",X"60",X"32",X"77",X"60",X"32",X"87",
		X"65",X"32",X"9A",X"65",X"32",X"9B",X"65",X"32",X"59",X"61",X"32",X"CF",X"61",X"32",X"E0",X"61",
		X"32",X"E1",X"61",X"3E",X"01",X"32",X"ED",X"61",X"CD",X"4D",X"2C",X"21",X"1A",X"90",X"11",X"20",
		X"00",X"3E",X"F0",X"06",X"20",X"77",X"E5",X"F5",X"7C",X"C6",X"08",X"67",X"3E",X"04",X"77",X"F1",
		X"E1",X"19",X"10",X"F1",X"CD",X"D7",X"38",X"3E",X"01",X"32",X"54",X"60",X"11",X"80",X"65",X"21",
		X"EE",X"38",X"01",X"04",X"00",X"ED",X"B0",X"11",X"9C",X"65",X"21",X"F2",X"38",X"01",X"04",X"00",
		X"ED",X"B0",X"3A",X"74",X"62",X"FE",X"01",X"CA",X"00",X"38",X"11",X"00",X"4C",X"21",X"86",X"92",
		X"3E",X"16",X"08",X"CD",X"F0",X"55",X"11",X"0B",X"4C",X"21",X"87",X"92",X"3E",X"16",X"08",X"CD",
		X"F0",X"55",X"11",X"16",X"4C",X"21",X"88",X"92",X"3E",X"16",X"08",X"CD",X"F0",X"55",X"11",X"21",
		X"4C",X"21",X"6B",X"92",X"3E",X"13",X"08",X"CD",X"F0",X"55",X"3A",X"00",X"B0",X"E6",X"20",X"FE",
		X"20",X"20",X"0A",X"3E",X"E1",X"32",X"8B",X"91",X"3E",X"13",X"32",X"8B",X"99",X"11",X"2A",X"4C",
		X"21",X"8E",X"93",X"3E",X"17",X"08",X"CD",X"F0",X"55",X"11",X"45",X"4C",X"21",X"8F",X"93",X"3E",
		X"17",X"08",X"CD",X"F0",X"55",X"11",X"60",X"4C",X"21",X"90",X"93",X"3E",X"17",X"08",X"CD",X"F0",
		X"55",X"11",X"7B",X"4C",X"21",X"52",X"92",X"3E",X"12",X"08",X"CD",X"F0",X"55",X"ED",X"56",X"FF",
		X"3A",X"26",X"60",X"F6",X"08",X"FB",X"32",X"26",X"60",X"3E",X"01",X"32",X"C7",X"61",X"CD",X"D7",
		X"38",X"3A",X"74",X"62",X"FE",X"01",X"28",X"08",X"3E",X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",
		X"3A",X"82",X"65",X"FE",X"20",X"20",X"D9",X"3A",X"26",X"60",X"F6",X"10",X"32",X"26",X"60",X"CD",
		X"D7",X"38",X"3A",X"82",X"65",X"FE",X"20",X"20",X"EE",X"11",X"94",X"65",X"21",X"F6",X"38",X"01",
		X"04",X"00",X"ED",X"B0",X"3A",X"26",X"60",X"F6",X"10",X"32",X"26",X"60",X"3E",X"80",X"32",X"27",
		X"60",X"CD",X"D7",X"38",X"3A",X"82",X"65",X"FE",X"F0",X"20",X"E9",X"CD",X"D7",X"38",X"3A",X"96",
		X"65",X"FE",X"D0",X"20",X"F6",X"3E",X"00",X"32",X"C7",X"61",X"3E",X"01",X"32",X"CF",X"61",X"3E",
		X"37",X"32",X"9C",X"65",X"3A",X"26",X"60",X"F6",X"08",X"32",X"26",X"60",X"3E",X"40",X"32",X"27",
		X"60",X"CD",X"D7",X"38",X"3A",X"82",X"65",X"FE",X"10",X"38",X"39",X"3A",X"74",X"62",X"FE",X"01",
		X"28",X"07",X"3A",X"48",X"92",X"FE",X"F6",X"20",X"2B",X"3A",X"82",X"65",X"FE",X"03",X"DD",X"21",
		X"94",X"65",X"FD",X"21",X"9C",X"65",X"0E",X"00",X"06",X"06",X"CD",X"D5",X"2A",X"FE",X"01",X"20",
		X"C3",X"CD",X"41",X"22",X"06",X"03",X"21",X"00",X"50",X"2B",X"CD",X"D7",X"38",X"7C",X"FE",X"00",
		X"20",X"F7",X"10",X"F2",X"3E",X"00",X"C3",X"69",X"5E",X"06",X"01",X"21",X"80",X"65",X"3E",X"00",
		X"32",X"54",X"60",X"CD",X"F1",X"29",X"C9",X"3A",X"00",X"60",X"FE",X"00",X"C8",X"3A",X"74",X"62",
		X"FE",X"01",X"C8",X"3E",X"00",X"32",X"ED",X"61",X"3A",X"00",X"B8",X"E1",X"18",X"D6",X"20",X"08",
		X"F0",X"C0",X"3A",X"28",X"E5",X"C0",X"31",X"0C",X"00",X"C0",X"CD",X"07",X"39",X"CD",X"24",X"39",
		X"CD",X"41",X"39",X"CD",X"5E",X"39",X"C9",X"3A",X"26",X"60",X"E6",X"01",X"47",X"3A",X"50",X"60",
		X"E6",X"01",X"B8",X"C8",X"3A",X"50",X"60",X"E6",X"01",X"FE",X"01",X"C0",X"3E",X"01",X"0E",X"01",
		X"CD",X"7B",X"39",X"C9",X"3A",X"26",X"60",X"E6",X"02",X"47",X"3A",X"50",X"60",X"E6",X"02",X"B8",
		X"C8",X"3A",X"50",X"60",X"E6",X"02",X"FE",X"02",X"C0",X"3E",X"02",X"0E",X"02",X"CD",X"7B",X"39",
		X"C9",X"3A",X"51",X"60",X"E6",X"01",X"47",X"3A",X"52",X"60",X"E6",X"01",X"B8",X"C8",X"3A",X"52",
		X"60",X"E6",X"01",X"FE",X"01",X"C0",X"3E",X"06",X"0E",X"05",X"CD",X"7B",X"39",X"C9",X"3A",X"51",
		X"60",X"E6",X"02",X"47",X"3A",X"52",X"60",X"E6",X"02",X"B8",X"C8",X"3A",X"52",X"60",X"E6",X"02",
		X"FE",X"02",X"C0",X"3E",X"0E",X"0E",X"0A",X"CD",X"7B",X"39",X"C9",X"F5",X"CD",X"F6",X"39",X"F1",
		X"47",X"3A",X"63",X"61",X"E6",X"04",X"FE",X"04",X"78",X"28",X"01",X"87",X"21",X"E4",X"61",X"86",
		X"77",X"FE",X"02",X"D4",X"97",X"39",X"C9",X"21",X"E4",X"61",X"7E",X"FE",X"02",X"D8",X"3A",X"00",
		X"60",X"FE",X"90",X"C8",X"C6",X"01",X"27",X"32",X"00",X"60",X"21",X"E4",X"61",X"35",X"35",X"21",
		X"68",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"CD",X"BE",X"39",X"18",X"D9",X"3A",X"00",
		X"60",X"E6",X"0F",X"32",X"9F",X"90",X"3A",X"00",X"60",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",
		X"0F",X"E6",X"0F",X"32",X"BF",X"90",X"3E",X"E0",X"06",X"07",X"21",X"9F",X"93",X"CD",X"BC",X"29",
		X"3A",X"56",X"60",X"FE",X"00",X"C8",X"21",X"9F",X"93",X"47",X"3E",X"CA",X"CD",X"BC",X"29",X"C9",
		X"01",X"01",X"01",X"00",X"01",X"00",X"79",X"21",X"E5",X"61",X"86",X"77",X"C9",X"3A",X"26",X"60",
		X"32",X"50",X"60",X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"38",X"D3",X"09",X"3E",
		X"0E",X"D3",X"08",X"DB",X"0C",X"2F",X"CD",X"3F",X"3A",X"CD",X"54",X"3A",X"32",X"26",X"60",X"3A",
		X"51",X"60",X"32",X"52",X"60",X"3E",X"0F",X"D3",X"08",X"DB",X"0C",X"2F",X"CD",X"3F",X"3A",X"32",
		X"51",X"60",X"3A",X"00",X"B0",X"2F",X"32",X"63",X"61",X"3E",X"01",X"32",X"07",X"A0",X"C9",X"F5",
		X"3A",X"ED",X"61",X"FE",X"01",X"28",X"09",X"3A",X"F2",X"61",X"FE",X"01",X"28",X"02",X"F1",X"C9",
		X"F1",X"E6",X"07",X"C9",X"47",X"3A",X"00",X"B0",X"2F",X"CB",X"07",X"E6",X"01",X"4F",X"3A",X"7C",
		X"61",X"A1",X"32",X"FD",X"61",X"FE",X"01",X"28",X"02",X"78",X"C9",X"3A",X"51",X"60",X"E6",X"F8",
		X"4F",X"78",X"E6",X"07",X"B1",X"C9",X"30",X"40",X"00",X"4C",X"A0",X"4E",X"21",X"47",X"00",X"45",
		X"02",X"4C",X"04",X"49",X"30",X"47",X"20",X"7F",X"30",X"6E",X"11",X"67",X"30",X"6D",X"10",X"C6",
		X"00",X"7D",X"84",X"4B",X"A1",X"CD",X"10",X"49",X"00",X"6D",X"00",X"4D",X"14",X"56",X"10",X"46",
		X"00",X"50",X"19",X"59",X"20",X"4A",X"20",X"4D",X"20",X"40",X"B1",X"42",X"00",X"64",X"10",X"49",
		X"04",X"59",X"24",X"60",X"20",X"4A",X"20",X"44",X"80",X"49",X"04",X"45",X"10",X"4D",X"00",X"4D",
		X"31",X"4B",X"02",X"4F",X"00",X"44",X"20",X"49",X"20",X"49",X"05",X"4C",X"23",X"CA",X"24",X"47",
		X"20",X"4A",X"00",X"41",X"81",X"FE",X"20",X"4E",X"10",X"6C",X"10",X"49",X"30",X"C4",X"20",X"4B",
		X"30",X"4B",X"21",X"69",X"10",X"4E",X"84",X"4C",X"04",X"46",X"82",X"43",X"B0",X"44",X"10",X"4D",
		X"00",X"41",X"10",X"45",X"B4",X"42",X"90",X"4C",X"06",X"40",X"21",X"67",X"02",X"CE",X"00",X"4C",
		X"CD",X"8C",X"3B",X"79",X"FE",X"00",X"C8",X"01",X"C7",X"61",X"D9",X"FD",X"21",X"C4",X"61",X"3E",
		X"3A",X"FD",X"77",X"04",X"3E",X"28",X"FD",X"77",X"05",X"3E",X"EC",X"32",X"CA",X"61",X"FD",X"56",
		X"01",X"FD",X"5E",X"00",X"CD",X"76",X"21",X"21",X"1B",X"3F",X"CD",X"18",X"20",X"3A",X"56",X"60",
		X"3C",X"32",X"56",X"60",X"3A",X"26",X"60",X"F6",X"10",X"32",X"26",X"60",X"AF",X"32",X"96",X"65",
		X"32",X"9A",X"65",X"3E",X"01",X"32",X"00",X"A0",X"32",X"F2",X"61",X"FB",X"CD",X"53",X"16",X"3A",
		X"82",X"65",X"FE",X"F0",X"20",X"DE",X"AF",X"32",X"F2",X"61",X"32",X"C7",X"61",X"F3",X"06",X"40",
		X"21",X"80",X"65",X"3E",X"00",X"77",X"23",X"10",X"FC",X"21",X"00",X"52",X"22",X"40",X"61",X"AF",
		X"32",X"42",X"61",X"3E",X"01",X"32",X"74",X"62",X"CD",X"00",X"37",X"AF",X"32",X"74",X"62",X"3C",
		X"32",X"54",X"60",X"CD",X"4F",X"35",X"31",X"F0",X"67",X"C3",X"2B",X"12",X"0E",X"00",X"FD",X"21",
		X"9C",X"60",X"06",X"36",X"FD",X"7E",X"00",X"FE",X"00",X"C0",X"FD",X"23",X"10",X"F6",X"C3",X"60",
		X"5E",X"21",X"F4",X"61",X"7E",X"47",X"3A",X"E8",X"61",X"B8",X"C8",X"FE",X"05",X"D0",X"21",X"94",
		X"5B",X"22",X"40",X"61",X"32",X"F4",X"61",X"AF",X"32",X"42",X"61",X"C9",X"3A",X"0D",X"60",X"32",
		X"98",X"60",X"FD",X"21",X"61",X"61",X"DD",X"21",X"84",X"65",X"CD",X"8C",X"55",X"3A",X"0D",X"60",
		X"FE",X"01",X"C8",X"DD",X"7E",X"03",X"FE",X"11",X"D8",X"3A",X"0D",X"60",X"FE",X"02",X"20",X"0D",
		X"11",X"DE",X"4B",X"AF",X"ED",X"5A",X"11",X"62",X"91",X"06",X"0F",X"18",X"0B",X"11",X"DE",X"47",
		X"AF",X"ED",X"5A",X"11",X"02",X"93",X"06",X"17",X"3E",X"FB",X"E5",X"AF",X"ED",X"52",X"E1",X"28",
		X"09",X"3E",X"FB",X"CD",X"2C",X"3C",X"13",X"10",X"EF",X"C9",X"DD",X"7E",X"03",X"E6",X"07",X"47",
		X"3E",X"F3",X"80",X"CD",X"2C",X"3C",X"06",X"03",X"13",X"C5",X"1A",X"01",X"08",X"00",X"21",X"3F",
		X"3C",X"ED",X"B1",X"3E",X"F3",X"CC",X"2C",X"3C",X"C1",X"10",X"ED",X"C9",X"12",X"C5",X"47",X"1A",
		X"B8",X"78",X"C1",X"20",X"F7",X"D5",X"7A",X"C6",X"08",X"57",X"3E",X"20",X"12",X"D1",X"C9",X"FB",
		X"FA",X"F9",X"F8",X"F7",X"F6",X"F5",X"F4",X"2A",X"91",X"60",X"22",X"FF",X"61",X"2A",X"93",X"60",
		X"22",X"01",X"62",X"2A",X"95",X"60",X"22",X"03",X"62",X"3A",X"0B",X"60",X"32",X"05",X"62",X"3A",
		X"98",X"60",X"32",X"F9",X"61",X"C9",X"2A",X"FF",X"61",X"22",X"91",X"60",X"2A",X"01",X"62",X"22",
		X"93",X"60",X"2A",X"03",X"62",X"22",X"95",X"60",X"3A",X"05",X"62",X"32",X"0B",X"60",X"3A",X"F9",
		X"61",X"32",X"98",X"60",X"C9",X"F5",X"D5",X"E5",X"06",X"00",X"CD",X"AA",X"3C",X"20",X"17",X"23",
		X"CD",X"AA",X"3C",X"20",X"11",X"11",X"1F",X"00",X"19",X"CD",X"AA",X"3C",X"20",X"08",X"23",X"CD",
		X"AA",X"3C",X"20",X"02",X"06",X"01",X"E1",X"D1",X"F1",X"C9",X"7E",X"FE",X"E0",X"C8",X"FE",X"49",
		X"C8",X"FE",X"4A",X"C8",X"FE",X"4B",X"C9",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"E1",X"C9",
		X"DD",X"21",X"CC",X"61",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"03",X"3E",X"FF",
		X"32",X"9F",X"65",X"C9",X"CD",X"75",X"55",X"CD",X"7A",X"3D",X"28",X"12",X"AF",X"32",X"77",X"60",
		X"3A",X"09",X"62",X"FE",X"01",X"20",X"07",X"CD",X"7C",X"22",X"AF",X"32",X"09",X"62",X"DD",X"21",
		X"8F",X"60",X"FD",X"21",X"57",X"61",X"21",X"98",X"65",X"22",X"15",X"62",X"2A",X"78",X"60",X"11",
		X"7B",X"60",X"3A",X"9A",X"60",X"32",X"98",X"60",X"01",X"12",X"62",X"CD",X"49",X"3D",X"CD",X"68",
		X"55",X"CD",X"7A",X"3D",X"28",X"12",X"AF",X"32",X"37",X"60",X"3A",X"08",X"62",X"FE",X"01",X"20",
		X"07",X"CD",X"41",X"22",X"AF",X"32",X"08",X"62",X"DD",X"21",X"4F",X"60",X"FD",X"21",X"56",X"61",
		X"21",X"94",X"65",X"22",X"15",X"62",X"2A",X"38",X"60",X"11",X"3B",X"60",X"3A",X"99",X"60",X"32",
		X"98",X"60",X"01",X"11",X"62",X"CD",X"49",X"3D",X"C9",X"DD",X"7E",X"00",X"FE",X"12",X"38",X"0E",
		X"CD",X"7A",X"3D",X"20",X"63",X"1A",X"FE",X"01",X"28",X"5E",X"3E",X"01",X"02",X"C9",X"0A",X"FE",
		X"01",X"28",X"5B",X"AF",X"C9",X"7E",X"E5",X"C5",X"01",X"02",X"00",X"21",X"78",X"3D",X"ED",X"B1",
		X"C1",X"E1",X"C8",X"AF",X"32",X"08",X"60",X"C9",X"E0",X"FB",X"7E",X"E5",X"C5",X"01",X"30",X"00",
		X"21",X"88",X"3D",X"ED",X"B1",X"C1",X"E1",X"C9",X"FF",X"FE",X"FD",X"FC",X"FB",X"FA",X"F9",X"E2",
		X"E1",X"E0",X"DF",X"DE",X"CF",X"CE",X"CA",X"BA",X"B7",X"A4",X"9B",X"9A",X"98",X"97",X"87",X"86",
		X"7E",X"7D",X"73",X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"68",X"67",X"66",X"64",X"63",X"62",X"5E",
		X"5D",X"52",X"45",X"44",X"41",X"3D",X"3C",X"29",X"2A",X"15",X"62",X"3E",X"22",X"77",X"AF",X"02",
		X"3E",X"01",X"FD",X"77",X"00",X"EB",X"11",X"04",X"00",X"AF",X"ED",X"52",X"77",X"21",X"37",X"04",
		X"22",X"54",X"61",X"AF",X"32",X"F5",X"61",X"3A",X"98",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"C0",
		X"21",X"4B",X"3F",X"CD",X"18",X"20",X"AF",X"32",X"53",X"61",X"C9",X"DD",X"E5",X"DD",X"2A",X"40",
		X"61",X"DD",X"7E",X"03",X"DD",X"E1",X"FE",X"FF",X"C9",X"3A",X"00",X"B8",X"DD",X"21",X"80",X"65",
		X"FD",X"21",X"A8",X"65",X"CD",X"01",X"10",X"DD",X"21",X"84",X"65",X"FD",X"21",X"A4",X"65",X"CD",
		X"01",X"10",X"DD",X"21",X"88",X"65",X"FD",X"21",X"AC",X"65",X"CD",X"01",X"10",X"DD",X"21",X"8C",
		X"65",X"FD",X"21",X"B0",X"65",X"CD",X"01",X"10",X"DD",X"21",X"90",X"65",X"FD",X"21",X"B4",X"65",
		X"CD",X"01",X"10",X"DD",X"21",X"9C",X"65",X"FD",X"21",X"A0",X"65",X"CD",X"01",X"10",X"AF",X"32",
		X"5F",X"98",X"3A",X"00",X"B0",X"2F",X"E6",X"80",X"CB",X"07",X"06",X"01",X"FE",X"00",X"28",X"07",
		X"47",X"3A",X"7C",X"61",X"2F",X"A0",X"47",X"48",X"06",X"08",X"11",X"04",X"00",X"21",X"A3",X"65",
		X"7E",X"FE",X"00",X"28",X"02",X"81",X"77",X"19",X"10",X"F6",X"21",X"AF",X"65",X"06",X"03",X"35",
		X"19",X"10",X"FC",X"79",X"FE",X"00",X"20",X"16",X"3A",X"0D",X"60",X"FE",X"01",X"28",X"0F",X"3A",
		X"ED",X"61",X"FE",X"01",X"28",X"08",X"3A",X"A6",X"65",X"3C",X"3C",X"32",X"A6",X"65",X"C9",X"00",
		X"00",X"B2",X"05",X"61",X"05",X"14",X"05",X"CC",X"04",X"86",X"04",X"45",X"04",X"08",X"04",X"CE",
		X"03",X"97",X"03",X"63",X"03",X"34",X"03",X"05",X"03",X"D9",X"02",X"B0",X"02",X"8A",X"02",X"66",
		X"02",X"43",X"02",X"22",X"02",X"04",X"02",X"E7",X"01",X"CB",X"01",X"B2",X"01",X"99",X"01",X"82",
		X"01",X"6D",X"01",X"58",X"01",X"45",X"01",X"33",X"01",X"22",X"01",X"11",X"01",X"02",X"01",X"F4",
		X"00",X"E6",X"00",X"D9",X"00",X"CD",X"00",X"C1",X"00",X"B6",X"00",X"AC",X"00",X"A2",X"00",X"9A",
		X"00",X"91",X"00",X"89",X"00",X"81",X"00",X"7A",X"00",X"73",X"00",X"6C",X"00",X"66",X"00",X"61",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"01",X"00",
		X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",
		X"01",X"46",X"24",X"4F",X"20",X"5C",X"14",X"4F",X"08",X"4F",X"21",X"47",X"19",X"43",X"00",X"46",
		X"84",X"43",X"13",X"46",X"34",X"4D",X"02",X"C0",X"00",X"65",X"90",X"46",X"20",X"44",X"00",X"4C",
		X"10",X"45",X"01",X"44",X"10",X"67",X"02",X"4E",X"00",X"4F",X"20",X"5C",X"00",X"49",X"00",X"44",
		X"00",X"48",X"0A",X"5C",X"20",X"49",X"00",X"4D",X"A0",X"40",X"A1",X"6A",X"A1",X"60",X"00",X"4C",
		X"00",X"4C",X"10",X"6B",X"24",X"5C",X"03",X"4E",X"20",X"4F",X"22",X"49",X"FF",X"BA",X"EA",X"97",
		X"A3",X"CA",X"01",X"4F",X"13",X"4B",X"10",X"47",X"21",X"5D",X"00",X"4C",X"10",X"C7",X"24",X"49",
		X"00",X"47",X"34",X"C5",X"15",X"46",X"30",X"CC",X"20",X"49",X"20",X"40",X"7F",X"B4",X"EF",X"BF",
		X"32",X"4D",X"28",X"6D",X"A0",X"58",X"02",X"48",X"10",X"41",X"91",X"49",X"1D",X"41",X"20",X"5A",
		X"31",X"5F",X"00",X"05",X"10",X"CF",X"30",X"48",X"0A",X"52",X"00",X"49",X"FD",X"B1",X"FF",X"B2",
		X"00",X"4F",X"09",X"6A",X"A0",X"4C",X"22",X"42",X"81",X"6D",X"02",X"42",X"31",X"4F",X"34",X"C4",
		X"80",X"47",X"00",X"42",X"10",X"41",X"10",X"4E",X"01",X"4D",X"00",X"41",X"FE",X"B5",X"CF",X"01",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"E0",
		X"02",X"E0",X"E0",X"E0",X"DB",X"71",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"A5",X"D8",X"B9",X"DB",X"DB",X"46",X"E0",X"E0",X"D7",X"E0",
		X"E0",X"00",X"E0",X"E0",X"DB",X"A5",X"D8",X"0B",X"E0",X"E0",X"CB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"46",X"4A",X"E0",X"DB",X"DB",X"DB",X"A6",X"D8",X"D8",X"BE",X"DB",X"46",X"E0",X"E0",X"D6",X"E0",
		X"22",X"00",X"E0",X"E0",X"DB",X"D1",X"72",X"48",X"E0",X"E0",X"D3",X"85",X"DB",X"DB",X"DB",X"DB",
		X"46",X"4B",X"49",X"DB",X"DB",X"DB",X"DB",X"BC",X"E0",X"E0",X"DB",X"46",X"4A",X"E0",X"D6",X"00",
		X"15",X"00",X"E0",X"DF",X"FB",X"FE",X"73",X"6E",X"DF",X"DF",X"6C",X"6A",X"86",X"E4",X"E4",X"E4",
		X"E4",X"E0",X"E0",X"E4",X"E4",X"E4",X"E4",X"6A",X"E0",X"E0",X"DB",X"46",X"4B",X"49",X"D6",X"00",
		X"29",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DC",X"E0",X"E0",X"D6",X"E0",
		X"11",X"00",X"E0",X"DE",X"FA",X"FD",X"74",X"6F",X"DE",X"DE",X"6D",X"6B",X"6B",X"87",X"E5",X"E5",
		X"E5",X"E5",X"E0",X"E0",X"E5",X"E5",X"E5",X"6B",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"D6",X"24",
		X"1C",X"00",X"E0",X"E0",X"DB",X"DB",X"75",X"48",X"E0",X"E0",X"D3",X"D8",X"D8",X"88",X"DB",X"DB",
		X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"48",X"4A",X"E0",X"DB",X"46",X"E0",X"E0",X"D6",X"19",
		X"20",X"E0",X"E0",X"E0",X"DB",X"DB",X"76",X"48",X"E0",X"E0",X"D3",X"D8",X"D8",X"89",X"DB",X"DB",
		X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"48",X"4B",X"49",X"DB",X"46",X"E0",X"E0",X"D6",X"14",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"AA",X"48",X"E0",X"E0",X"D3",X"D8",X"8A",X"E4",X"FE",X"FE",
		X"FE",X"F9",X"DF",X"DF",X"DB",X"DB",X"A7",X"48",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"D5",X"15",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"77",X"D8",X"48",X"4A",X"E0",X"D3",X"8B",X"DB",X"E0",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"DB",X"DB",X"A8",X"48",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"D4",X"22",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"78",X"D8",X"48",X"4B",X"49",X"C9",X"8C",X"DB",X"E0",X"DE",X"FA",
		X"FD",X"FC",X"DE",X"DE",X"DB",X"DB",X"A9",X"48",X"4A",X"E0",X"DB",X"46",X"E0",X"E0",X"D3",X"13",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"79",X"D8",X"48",X"E0",X"E0",X"C8",X"DB",X"DB",X"E0",X"E0",X"DB",
		X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"AA",X"48",X"4B",X"49",X"DB",X"46",X"E0",X"E0",X"D3",X"E0",
		X"23",X"00",X"E0",X"E0",X"DB",X"7A",X"D8",X"48",X"E0",X"E0",X"C7",X"DB",X"EA",X"E0",X"F7",X"DB",
		X"DB",X"DB",X"F0",X"E0",X"F1",X"9F",X"D8",X"48",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"D3",X"E0",
		X"25",X"00",X"E0",X"E0",X"DB",X"AA",X"D8",X"48",X"E0",X"E0",X"C6",X"DB",X"EB",X"E0",X"F6",X"DB",
		X"DB",X"DB",X"EF",X"E0",X"F2",X"A0",X"D8",X"48",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"D3",X"E0",
		X"1E",X"05",X"E0",X"E0",X"DB",X"D8",X"D8",X"48",X"E0",X"E0",X"C5",X"DB",X"EC",X"E0",X"F5",X"DB",
		X"DB",X"DB",X"EE",X"E0",X"F3",X"A1",X"D8",X"48",X"E0",X"E0",X"DB",X"47",X"E0",X"E0",X"D3",X"E0",
		X"1F",X"09",X"E0",X"E0",X"DB",X"D8",X"D8",X"0B",X"E0",X"E0",X"C4",X"DB",X"ED",X"E0",X"F4",X"DB",
		X"DB",X"DB",X"ED",X"E0",X"F4",X"AA",X"D8",X"48",X"E0",X"E0",X"C5",X"48",X"E0",X"E0",X"D3",X"E0",
		X"12",X"E0",X"E0",X"E0",X"DB",X"AD",X"D8",X"48",X"E0",X"E0",X"C3",X"DB",X"EE",X"E0",X"F3",X"DB",
		X"DB",X"DB",X"EC",X"E0",X"F5",X"D8",X"D8",X"48",X"E0",X"E0",X"C6",X"48",X"E0",X"E0",X"D2",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"AE",X"D8",X"48",X"4A",X"E0",X"C2",X"DB",X"EF",X"E0",X"F2",X"DB",
		X"DB",X"DB",X"EB",X"E0",X"F6",X"D8",X"D8",X"48",X"4A",X"E0",X"C7",X"0B",X"E0",X"E0",X"D1",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"7B",X"D8",X"48",X"4B",X"49",X"C1",X"DB",X"F0",X"E0",X"F1",X"DB",
		X"DB",X"DB",X"EA",X"E0",X"F7",X"A2",X"D8",X"48",X"4B",X"49",X"C8",X"48",X"4A",X"E0",X"D0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"7C",X"D8",X"48",X"E0",X"E0",X"C0",X"96",X"E0",X"E0",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"E0",X"E0",X"A3",X"D8",X"48",X"E0",X"E0",X"C9",X"48",X"4B",X"49",X"CD",X"E0",
		X"01",X"E0",X"E0",X"DF",X"FB",X"7D",X"68",X"6E",X"DF",X"DF",X"6C",X"97",X"DF",X"DF",X"FB",X"FE",
		X"FE",X"FE",X"F9",X"DF",X"DF",X"A4",X"68",X"B7",X"DF",X"DF",X"FB",X"CE",X"DF",X"DF",X"D3",X"E0",
		X"E0",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D3",X"E0",
		X"22",X"00",X"E0",X"DE",X"FA",X"FD",X"7E",X"67",X"67",X"67",X"67",X"67",X"98",X"FC",X"DE",X"DE",
		X"FA",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"BA",X"FD",X"FD",X"CF",X"DE",X"DE",X"D3",X"E0",
		X"15",X"00",X"E0",X"E0",X"DB",X"DB",X"DB",X"7F",X"D8",X"D8",X"D8",X"D8",X"99",X"DB",X"E0",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"BB",X"DB",X"DB",X"46",X"4A",X"E0",X"D3",X"E0",
		X"29",X"00",X"E0",X"E0",X"DB",X"DB",X"DB",X"80",X"D8",X"D8",X"48",X"6A",X"9A",X"F9",X"DF",X"DF",
		X"FB",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"D8",X"BF",X"DB",X"46",X"4B",X"49",X"D3",X"E0",
		X"11",X"00",X"E0",X"E0",X"DB",X"DB",X"DB",X"81",X"D8",X"D8",X"48",X"E0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D8",X"C0",X"C1",X"46",X"E0",X"E0",X"D3",X"E0",
		X"1C",X"00",X"E0",X"E0",X"DB",X"DB",X"DB",X"82",X"D8",X"D8",X"48",X"6B",X"9B",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"70",X"BC",X"D8",X"C2",X"C3",X"DB",X"DB",X"DA",X"E0",
		X"20",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"83",X"D8",X"D8",X"D8",X"91",X"9C",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"BD",X"D8",X"D8",X"C4",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"02",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"5F",X"BC",X"D8",X"D8",X"5C",X"DB",X"DB",X"DB",X"51",
		X"48",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"3E",X"48",X"E0",X"E0",X"C4",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"46",X"E0",X"DF",X"FB",X"5E",X"68",X"68",X"5D",X"F9",X"52",X"52",X"DB",
		X"32",X"E0",X"E0",X"32",X"DB",X"DB",X"DB",X"59",X"48",X"E0",X"E0",X"B8",X"DB",X"DB",X"DB",X"E0",
		X"22",X"E0",X"E0",X"E0",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",
		X"46",X"E0",X"E0",X"33",X"DB",X"DB",X"DB",X"3F",X"0B",X"E0",X"E0",X"B9",X"E0",X"E0",X"D6",X"E0",
		X"15",X"E0",X"E0",X"E0",X"46",X"E0",X"DE",X"FA",X"67",X"67",X"67",X"63",X"FC",X"DE",X"DE",X"DB",
		X"46",X"E0",X"E0",X"D8",X"31",X"DB",X"DB",X"5F",X"48",X"E0",X"E0",X"C1",X"E0",X"E0",X"D6",X"E0",
		X"29",X"E0",X"E0",X"E0",X"46",X"4A",X"E0",X"60",X"D8",X"D8",X"E0",X"E0",X"DB",X"E0",X"E0",X"DB",
		X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"D6",X"E0",
		X"11",X"E0",X"E0",X"E0",X"46",X"4B",X"49",X"61",X"D8",X"D8",X"E0",X"E0",X"DB",X"E0",X"E0",X"DB",
		X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"DF",X"DF",X"DF",X"6C",X"DF",X"DF",X"D6",X"24",
		X"1C",X"E0",X"E0",X"E0",X"46",X"E0",X"DF",X"62",X"68",X"6E",X"DF",X"DF",X"DB",X"E0",X"E0",X"DB",
		X"46",X"E0",X"E0",X"D8",X"D8",X"34",X"EA",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"19",
		X"20",X"E0",X"E0",X"E0",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",X"E0",X"E0",X"DB",
		X"46",X"4A",X"E0",X"48",X"D8",X"35",X"EA",X"E0",X"DE",X"FA",X"41",X"6F",X"DE",X"DE",X"D6",X"14",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"5A",X"67",X"67",X"67",X"67",X"64",X"FD",X"DB",X"E0",X"E0",X"DB",
		X"46",X"4B",X"49",X"30",X"D8",X"4D",X"EA",X"E0",X"F7",X"DB",X"80",X"48",X"4A",X"E0",X"D6",X"15",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"C9",X"D8",X"36",X"EB",X"E0",X"F6",X"DB",X"42",X"48",X"4B",X"49",X"BF",X"22",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"82",X"D8",X"D8",X"EC",X"E0",X"F5",X"DB",X"DB",X"48",X"E0",X"E0",X"BE",X"13",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"AA",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"46",X"E0",X"E0",X"C6",X"D8",X"37",X"ED",X"E0",X"F4",X"DB",X"DB",X"48",X"E0",X"E0",X"BD",X"E0",
		X"23",X"E0",X"E0",X"E0",X"DB",X"D8",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"46",X"4A",X"E0",X"C7",X"D8",X"38",X"EE",X"E0",X"F3",X"DB",X"C5",X"48",X"E0",X"E0",X"BC",X"E0",
		X"25",X"E0",X"E0",X"E0",X"DB",X"D8",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"46",X"4B",X"49",X"76",X"D8",X"39",X"EF",X"E0",X"F2",X"DB",X"CC",X"0B",X"E0",X"E0",X"D6",X"E0",
		X"1E",X"E0",X"E0",X"E0",X"DB",X"AD",X"D8",X"0B",X"E0",X"E0",X"CB",X"46",X"DB",X"DB",X"DB",X"DB",
		X"46",X"E0",X"E0",X"AA",X"D8",X"3A",X"F0",X"E0",X"F1",X"DB",X"CD",X"48",X"4A",X"E0",X"D6",X"E0",
		X"1F",X"E0",X"E0",X"E0",X"DB",X"AE",X"D8",X"48",X"4A",X"E0",X"D3",X"40",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"E0",X"D8",X"D8",X"3B",X"E0",X"E0",X"DB",X"C5",X"D8",X"48",X"4B",X"49",X"D6",X"E0",
		X"12",X"E0",X"E0",X"E0",X"DB",X"7B",X"D8",X"48",X"4B",X"49",X"D3",X"48",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"DF",X"6C",X"68",X"3C",X"DF",X"DF",X"FB",X"44",X"68",X"6E",X"DF",X"DF",X"D6",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"7C",X"D8",X"48",X"E0",X"E0",X"D3",X"48",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"D1",X"D8",X"48",X"E0",X"E0",X"D3",X"48",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"DE",X"6D",X"67",X"3D",X"FD",X"FC",X"E0",X"E0",X"6D",X"6F",X"DE",X"DE",X"D6",X"E0",
		X"E0",X"E0",X"E0",X"DF",X"FB",X"FE",X"5E",X"6E",X"DF",X"DF",X"D3",X"48",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"E0",X"A2",X"D8",X"92",X"DB",X"DB",X"E0",X"E0",X"D8",X"48",X"E0",X"E0",X"D6",X"E0",
		X"01",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D3",X"48",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"E0",X"A3",X"D8",X"93",X"DB",X"DB",X"E0",X"E0",X"D8",X"48",X"E0",X"E0",X"D6",X"E0",
		X"E0",X"E0",X"E0",X"DE",X"FA",X"FD",X"67",X"6F",X"DE",X"DE",X"D3",X"48",X"4A",X"E0",X"DB",X"DB",
		X"46",X"E0",X"E0",X"59",X"D8",X"4F",X"DB",X"DB",X"E0",X"E0",X"D8",X"48",X"4A",X"E0",X"D6",X"E0",
		X"22",X"E0",X"E0",X"E0",X"DB",X"77",X"D8",X"48",X"4A",X"E0",X"D3",X"3F",X"4B",X"49",X"DB",X"DB",
		X"46",X"E0",X"E0",X"58",X"D8",X"4D",X"DB",X"DB",X"0A",X"09",X"57",X"48",X"4B",X"49",X"D6",X"E0",
		X"15",X"E0",X"E0",X"E0",X"DB",X"78",X"D8",X"48",X"4B",X"49",X"C9",X"3E",X"E0",X"E0",X"DB",X"DB",
		X"46",X"E0",X"E0",X"5F",X"72",X"D8",X"E0",X"E0",X"E0",X"E0",X"48",X"48",X"E0",X"E0",X"D6",X"E0",
		X"29",X"E0",X"E0",X"E0",X"DB",X"79",X"D8",X"48",X"E0",X"DF",X"66",X"F9",X"DF",X"DF",X"DB",X"DB",
		X"46",X"E0",X"E0",X"DB",X"56",X"D8",X"E0",X"E0",X"E0",X"E0",X"A5",X"48",X"E0",X"E0",X"BB",X"E0",
		X"11",X"E0",X"E0",X"E0",X"DB",X"7A",X"D8",X"48",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",X"DB",
		X"46",X"E0",X"E0",X"DB",X"55",X"D8",X"E0",X"E0",X"E0",X"E0",X"49",X"35",X"E0",X"E0",X"D3",X"E0",
		X"1C",X"E0",X"E0",X"E0",X"DB",X"AA",X"D8",X"48",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"DB",X"DB",
		X"46",X"4A",X"E0",X"DB",X"DB",X"54",X"E0",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"D3",X"E0",
		X"20",X"E0",X"E0",X"E0",X"C5",X"D8",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"46",X"4B",X"49",X"DB",X"DB",X"53",X"D8",X"C0",X"C1",X"DB",X"DB",X"46",X"E0",X"E0",X"D3",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"02",X"E0",X"E0",X"E0",X"46",X"83",X"D8",X"D8",X"D8",X"0F",X"DB",X"DB",X"DB",X"DB",X"A8",X"D8",
		X"D8",X"AB",X"21",X"77",X"D8",X"D8",X"D8",X"D8",X"D8",X"8B",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"46",X"10",X"68",X"68",X"68",X"9A",X"FE",X"DB",X"DB",X"DB",X"11",X"D8",
		X"D8",X"48",X"E4",X"44",X"68",X"68",X"68",X"68",X"6E",X"23",X"52",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"22",X"E0",X"E0",X"E0",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",X"DB",X"DB",X"17",X"D8",
		X"D8",X"48",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"15",X"E0",X"E0",X"E0",X"46",X"E0",X"DE",X"6D",X"6F",X"DE",X"DE",X"DB",X"DB",X"A7",X"D8",X"D8",
		X"D8",X"48",X"E0",X"DE",X"6D",X"67",X"67",X"67",X"24",X"DE",X"DE",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"29",X"E0",X"E0",X"DF",X"FB",X"DF",X"DF",X"D8",X"48",X"E0",X"DF",X"FB",X"FE",X"44",X"68",X"68",
		X"68",X"6E",X"DF",X"DF",X"D8",X"D8",X"D8",X"D8",X"36",X"4A",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"11",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"D8",X"48",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"D8",X"D8",X"D8",X"D8",X"37",X"4B",X"49",X"D6",X"DB",X"DB",X"DB",X"24",
		X"1C",X"E0",X"E0",X"DE",X"FA",X"DE",X"DE",X"D8",X"48",X"E0",X"DE",X"FA",X"FD",X"1B",X"67",X"67",
		X"67",X"6F",X"DE",X"DE",X"3E",X"D8",X"D8",X"D8",X"38",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"19",
		X"20",X"E0",X"E0",X"E0",X"46",X"4A",X"E0",X"D8",X"48",X"4A",X"E0",X"DB",X"DB",X"42",X"BC",X"D8",
		X"D8",X"48",X"E0",X"E0",X"7B",X"D8",X"D8",X"D8",X"39",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"14",
		X"E0",X"E0",X"E0",X"E0",X"46",X"4B",X"49",X"D8",X"48",X"4B",X"49",X"DB",X"DB",X"DB",X"50",X"D8",
		X"D8",X"48",X"E0",X"DF",X"22",X"68",X"68",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"15",
		X"E0",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"D8",X"48",X"E0",X"E0",X"96",X"DB",X"DB",X"51",X"1D",
		X"D8",X"48",X"E0",X"FF",X"FF",X"FF",X"FF",X"D8",X"48",X"4A",X"E0",X"D6",X"DB",X"DB",X"DB",X"22",
		X"E0",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"0E",X"48",X"E0",X"E0",X"16",X"DB",X"DB",X"DB",X"1C",
		X"D8",X"48",X"E0",X"DE",X"26",X"DE",X"DE",X"D8",X"48",X"4B",X"49",X"D6",X"DB",X"DB",X"DB",X"13",
		X"E0",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"0D",X"48",X"E0",X"E0",X"15",X"96",X"DB",X"DB",X"0C",
		X"68",X"6E",X"DF",X"DF",X"46",X"E0",X"DF",X"6C",X"6E",X"DF",X"DF",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"23",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"DB",X"34",X"4A",X"E0",X"D8",X"13",X"DB",X"DB",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"25",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"DB",X"33",X"4B",X"49",X"D8",X"14",X"31",X"DB",X"E0",
		X"E0",X"6D",X"67",X"27",X"46",X"E0",X"DE",X"25",X"6F",X"DE",X"DE",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"1E",X"E0",X"E0",X"E0",X"46",X"E0",X"DF",X"FB",X"29",X"DF",X"DF",X"D8",X"D8",X"12",X"EA",X"E0",
		X"F7",X"48",X"D8",X"35",X"46",X"4A",X"E0",X"80",X"48",X"4A",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"1F",X"E0",X"E0",X"E0",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"D8",X"D8",X"36",X"EB",X"E0",
		X"F6",X"30",X"D8",X"4D",X"46",X"4B",X"49",X"42",X"48",X"4B",X"49",X"BF",X"DB",X"DB",X"DB",X"E0",
		X"12",X"E0",X"E0",X"E0",X"46",X"E0",X"DE",X"FA",X"74",X"67",X"67",X"D8",X"D8",X"AB",X"EC",X"E0",
		X"F5",X"C9",X"D8",X"36",X"46",X"E0",X"E0",X"DB",X"3C",X"E0",X"E0",X"BE",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"DB",X"75",X"D8",X"D8",X"D8",X"D8",X"28",X"ED",X"E0",
		X"F4",X"82",X"D8",X"D8",X"46",X"E0",X"E0",X"DB",X"3D",X"E0",X"E0",X"BD",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"46",X"4A",X"E0",X"DB",X"76",X"D8",X"D8",X"D8",X"D8",X"2B",X"EE",X"E0",
		X"F3",X"C6",X"D8",X"37",X"46",X"E0",X"E0",X"C5",X"48",X"E0",X"E0",X"BC",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"46",X"4B",X"49",X"DB",X"AA",X"D8",X"D8",X"D8",X"8B",X"DB",X"EF",X"E0",
		X"F2",X"C7",X"D8",X"38",X"46",X"4A",X"E0",X"CC",X"0B",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"01",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"77",X"D8",X"D8",X"D8",X"D8",X"8C",X"DB",X"F0",X"E0",
		X"F1",X"76",X"D8",X"39",X"46",X"4B",X"49",X"CD",X"48",X"4A",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"78",X"D8",X"D8",X"D8",X"8E",X"DB",X"DB",X"E0",X"E0",
		X"F8",X"AA",X"D8",X"3A",X"46",X"E0",X"E0",X"B1",X"48",X"4B",X"49",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"22",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"15",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"29",X"E0",X"E0",X"E0",X"46",X"4A",X"E0",X"D8",X"D8",X"D8",X"D8",X"B4",X"DB",X"DB",X"DB",X"DB",
		X"3B",X"4A",X"E0",X"DB",X"DB",X"DB",X"59",X"D8",X"48",X"4A",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"11",X"E0",X"E0",X"E0",X"46",X"4B",X"49",X"D8",X"D8",X"D8",X"D8",X"2A",X"DB",X"DB",X"DB",X"DB",
		X"3A",X"4B",X"49",X"DB",X"DB",X"DB",X"C8",X"D8",X"48",X"4B",X"49",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"1C",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"AD",X"D8",X"D8",X"D8",X"92",X"DB",X"DB",X"DB",X"C5",
		X"48",X"E0",X"E0",X"DB",X"DB",X"DB",X"C9",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"20",X"E0",X"E0",X"E0",X"46",X"E0",X"E0",X"AE",X"D8",X"D8",X"D8",X"93",X"DB",X"DB",X"DB",X"42",
		X"48",X"E0",X"E0",X"DB",X"DB",X"DB",X"46",X"D8",X"48",X"E0",X"E0",X"D6",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"E0",X"E0",X"E0",X"E0",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"FF",X"FE",X"FD",X"FC",X"E5",X"E5",X"EE",X"ED",X"EC",X"E5",X"3F",X"FB",X"FA",X"F9",X"F8",X"F4",
		X"F2",X"F0",X"EB",X"EA",X"E9",X"3F",X"E5",X"F7",X"F6",X"F5",X"F3",X"F1",X"EF",X"E8",X"E7",X"E6",
		X"3F",X"E4",X"E3",X"E2",X"E1",X"E2",X"E0",X"DF",X"E2",X"3F",X"91",X"91",X"91",X"D9",X"D8",X"D7",
		X"91",X"D6",X"D5",X"91",X"D4",X"D3",X"D2",X"D1",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",
		X"C8",X"91",X"91",X"91",X"3F",X"91",X"91",X"91",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",
		X"BF",X"BE",X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"B7",X"B6",X"B5",X"B4",X"91",X"91",X"91",X"3F",
		X"91",X"91",X"91",X"B3",X"B2",X"B1",X"B0",X"AF",X"AE",X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",
		X"A6",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",X"9F",X"91",X"91",X"3F",X"DE",X"91",X"DD",X"DC",X"DB",
		X"DA",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8A",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"3F",X"8C",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"8D",X"3F",X"85",X"84",X"83",X"82",X"81",X"80",X"7F",X"91",X"91",X"3F",
		X"91",X"54",X"89",X"88",X"87",X"86",X"91",X"91",X"91",X"3F",X"7E",X"7D",X"7C",X"7B",X"7A",X"91",
		X"91",X"91",X"91",X"3F",X"79",X"78",X"77",X"76",X"75",X"74",X"91",X"91",X"91",X"3F",X"73",X"72",
		X"71",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"3F",X"91",X"91",X"6A",X"69",X"68",X"67",X"66",X"91",
		X"91",X"3F",X"91",X"65",X"64",X"63",X"62",X"91",X"91",X"91",X"91",X"3F",X"61",X"60",X"5F",X"5E",
		X"5D",X"91",X"91",X"91",X"91",X"3F",X"5A",X"59",X"91",X"58",X"57",X"3F",X"5C",X"3F",X"5B",X"3F",
		X"56",X"3F",X"55",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"14",X"08",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"1B",X"08",X"0A",
		X"00",X"1A",X"0F",X"0A",X"00",X"1B",X"00",X"0A",X"00",X"1A",X"00",X"0A",X"00",X"1B",X"00",X"0A",
		X"00",X"0F",X"08",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"1B",X"08",X"0A",
		X"00",X"1A",X"0F",X"0A",X"00",X"1B",X"00",X"0A",X"30",X"1A",X"00",X"0A",X"2E",X"1B",X"00",X"0A",
		X"2C",X"14",X"08",X"0A",X"00",X"00",X"00",X"0A",X"2C",X"00",X"00",X"0A",X"2E",X"1B",X"08",X"0A",
		X"2C",X"1A",X"0F",X"0A",X"00",X"1B",X"00",X"0A",X"24",X"1A",X"00",X"0A",X"25",X"1B",X"00",X"0A",
		X"27",X"14",X"08",X"0A",X"29",X"00",X"00",X"0A",X"27",X"00",X"00",X"0A",X"24",X"1B",X"08",X"0A",
		X"27",X"1A",X"0F",X"0A",X"00",X"1B",X"00",X"0A",X"2C",X"1A",X"00",X"0A",X"2E",X"1B",X"00",X"0A",
		X"30",X"14",X"08",X"0A",X"00",X"00",X"00",X"0A",X"30",X"00",X"00",X"0A",X"00",X"1B",X"08",X"0A",
		X"30",X"1A",X"0F",X"0A",X"2E",X"1B",X"00",X"0A",X"2C",X"1A",X"00",X"0A",X"2E",X"1B",X"00",X"0A",
		X"30",X"0F",X"03",X"0A",X"00",X"00",X"00",X"0A",X"2E",X"00",X"00",X"0A",X"00",X"00",X"03",X"0A",
		X"2E",X"0F",X"0A",X"0A",X"00",X"00",X"00",X"0A",X"30",X"1A",X"00",X"0A",X"2E",X"1B",X"00",X"0A",
		X"2C",X"14",X"08",X"0A",X"00",X"00",X"00",X"0A",X"2C",X"00",X"00",X"0A",X"2E",X"1B",X"08",X"0A",
		X"2C",X"1A",X"0F",X"0A",X"00",X"1B",X"00",X"0A",X"24",X"1A",X"00",X"0A",X"25",X"1B",X"00",X"0A",
		X"27",X"14",X"08",X"0A",X"29",X"00",X"00",X"0A",X"27",X"00",X"00",X"0A",X"24",X"1B",X"08",X"0A",
		X"27",X"1A",X"0F",X"0A",X"00",X"1B",X"00",X"0A",X"2C",X"1A",X"00",X"0A",X"2E",X"1B",X"00",X"0A",
		X"30",X"14",X"08",X"0A",X"00",X"00",X"00",X"0A",X"30",X"00",X"00",X"0A",X"00",X"1B",X"08",X"0A",
		X"30",X"1A",X"0F",X"0A",X"2E",X"1B",X"00",X"0A",X"2C",X"1A",X"00",X"0A",X"2E",X"1B",X"00",X"0A",
		X"30",X"0F",X"03",X"0A",X"00",X"00",X"00",X"0A",X"2E",X"13",X"07",X"0A",X"00",X"00",X"00",X"0A",
		X"2C",X"14",X"08",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"FF",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"0F",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",
		X"14",X"22",X"08",X"0A",X"00",X"24",X"00",X"0A",X"00",X"2C",X"00",X"0A",X"00",X"27",X"08",X"0A",
		X"14",X"22",X"03",X"0A",X"00",X"24",X"00",X"0A",X"00",X"2C",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"11",X"22",X"0C",X"0A",X"00",X"24",X"00",X"0A",X"0F",X"2C",X"00",X"0A",X"00",X"27",X"0C",X"0A",
		X"0F",X"22",X"03",X"0A",X"00",X"24",X"00",X"0A",X"11",X"1D",X"00",X"0A",X"00",X"1B",X"00",X"0A",
		X"14",X"20",X"08",X"0A",X"00",X"24",X"00",X"0A",X"00",X"27",X"00",X"0A",X"00",X"2C",X"08",X"0A",
		X"00",X"27",X"03",X"0A",X"00",X"20",X"00",X"0A",X"00",X"24",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"00",X"20",X"0C",X"0A",X"00",X"24",X"00",X"0A",X"00",X"27",X"00",X"0A",X"00",X"2C",X"0C",X"0A",
		X"14",X"27",X"03",X"0A",X"00",X"20",X"00",X"0A",X"16",X"24",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"18",X"22",X"08",X"0A",X"00",X"24",X"00",X"0A",X"00",X"2C",X"00",X"0A",X"00",X"27",X"08",X"0A",
		X"18",X"22",X"03",X"0A",X"00",X"24",X"00",X"0A",X"00",X"2C",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"1B",X"22",X"0C",X"0A",X"00",X"24",X"00",X"0A",X"18",X"2C",X"00",X"0A",X"00",X"27",X"0C",X"0A",
		X"16",X"22",X"03",X"0A",X"00",X"24",X"00",X"0A",X"14",X"1D",X"00",X"0A",X"00",X"1B",X"00",X"0A",
		X"16",X"22",X"0A",X"0A",X"00",X"27",X"00",X"0A",X"00",X"2B",X"00",X"0A",X"00",X"2C",X"0A",X"0A",
		X"00",X"2B",X"03",X"0A",X"00",X"27",X"00",X"0A",X"00",X"22",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"00",X"22",X"0D",X"0A",X"00",X"27",X"00",X"0A",X"00",X"2B",X"00",X"0A",X"00",X"2C",X"0D",X"0A",
		X"1B",X"2B",X"03",X"0A",X"00",X"27",X"00",X"0A",X"19",X"22",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"18",X"22",X"08",X"0A",X"00",X"24",X"00",X"0A",X"00",X"2C",X"00",X"0A",X"00",X"27",X"08",X"0A",
		X"18",X"22",X"03",X"0A",X"00",X"24",X"00",X"0A",X"00",X"2C",X"00",X"0A",X"00",X"27",X"00",X"0A",
		X"16",X"22",X"0C",X"0A",X"00",X"24",X"00",X"0A",X"14",X"2C",X"00",X"0A",X"00",X"27",X"0C",X"0A",
		X"14",X"22",X"03",X"0A",X"00",X"24",X"00",X"0A",X"12",X"1D",X"00",X"0A",X"00",X"1B",X"00",X"0A",
		X"11",X"1D",X"0D",X"0A",X"00",X"20",X"00",X"0A",X"00",X"25",X"00",X"0A",X"00",X"27",X"0D",X"0A",
		X"11",X"25",X"08",X"0A",X"00",X"22",X"00",X"0A",X"00",X"20",X"00",X"0A",X"00",X"1D",X"00",X"0A",
		X"16",X"1C",X"05",X"0A",X"00",X"20",X"00",X"0A",X"14",X"25",X"00",X"0A",X"00",X"27",X"05",X"0A",
		X"13",X"25",X"01",X"0A",X"00",X"22",X"00",X"0A",X"11",X"20",X"00",X"0A",X"00",X"1C",X"00",X"0A",
		X"0F",X"1B",X"08",X"0A",X"00",X"20",X"00",X"0A",X"00",X"24",X"00",X"0A",X"00",X"25",X"08",X"0A",
		X"0F",X"24",X"03",X"0A",X"00",X"22",X"00",X"0A",X"00",X"20",X"00",X"0A",X"00",X"1D",X"00",X"0A",
		X"18",X"1B",X"0A",X"0A",X"00",X"1F",X"00",X"0A",X"16",X"22",X"00",X"0A",X"00",X"24",X"0A",X"0A",
		X"14",X"22",X"03",X"0A",X"00",X"1F",X"00",X"0A",X"13",X"1B",X"00",X"0A",X"00",X"1F",X"00",X"0A",
		X"14",X"20",X"08",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"FF",X"0E",X"60",X"6F",X"37",X"78",X"DE",X"FB",X"92",X"9B",X"5E",X"7F",X"9E",
		X"5B",X"5C",X"FF",X"9A",X"9C",X"4A",X"FF",X"5E",X"FD",X"7E",X"BF",X"DF",X"5F",X"5E",X"FF",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"ED",X"61",X"FE",X"01",X"C8",X"3A",X"7C",X"61",X"FE",X"00",X"C2",X"31",X"55",X"DD",X"21",
		X"76",X"61",X"AF",X"7D",X"47",X"DD",X"7E",X"00",X"80",X"27",X"DD",X"77",X"00",X"7C",X"47",X"DD",
		X"7E",X"01",X"88",X"27",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"CE",X"00",X"27",X"DD",X"77",X"02",
		X"C9",X"DD",X"21",X"79",X"61",X"18",X"DB",X"FD",X"7E",X"02",X"47",X"DD",X"7E",X"02",X"CD",X"4E",
		X"55",X"FD",X"7E",X"03",X"47",X"DD",X"7E",X"03",X"CD",X"4E",X"55",X"3E",X"01",X"C9",X"4F",X"C6",
		X"0B",X"B8",X"38",X"07",X"79",X"D6",X"08",X"B8",X"30",X"01",X"C9",X"F1",X"AF",X"C9",X"DD",X"21",
		X"80",X"65",X"FD",X"21",X"09",X"60",X"18",X"1A",X"DD",X"21",X"94",X"65",X"FD",X"21",X"38",X"60",
		X"3A",X"99",X"60",X"18",X"10",X"DD",X"21",X"98",X"65",X"FD",X"21",X"78",X"60",X"3A",X"9A",X"60",
		X"18",X"03",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",X"8C",X"55",X"C9",X"CD",X"AC",X"55",X"CD",
		X"9A",X"55",X"FD",X"75",X"00",X"FD",X"74",X"01",X"C9",X"C9",X"DD",X"7E",X"03",X"C6",X"10",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"C9",X"DD",X"7E",X"02",X"C6",
		X"07",X"2F",X"CB",X"3F",X"C3",X"CD",X"5B",X"00",X"47",X"11",X"20",X"00",X"21",X"00",X"40",X"19",
		X"10",X"FD",X"3A",X"98",X"60",X"FE",X"01",X"C8",X"FE",X"02",X"20",X"05",X"7C",X"C6",X"04",X"67",
		X"C9",X"FE",X"03",X"C0",X"7C",X"C6",X"08",X"67",X"C9",X"01",X"E0",X"FF",X"1A",X"FE",X"3F",X"C8",
		X"D6",X"30",X"77",X"E5",X"7C",X"C6",X"08",X"67",X"3E",X"00",X"77",X"E1",X"13",X"09",X"18",X"E9",
		X"01",X"E0",X"FF",X"1A",X"FE",X"3F",X"C8",X"77",X"E5",X"7C",X"C6",X"08",X"67",X"08",X"77",X"08",
		X"E1",X"13",X"09",X"18",X"EB",X"11",X"20",X"00",X"06",X"1C",X"77",X"19",X"10",X"FC",X"C9",X"DD",
		X"21",X"76",X"61",X"21",X"E1",X"92",X"CD",X"3C",X"56",X"DD",X"21",X"79",X"61",X"21",X"61",X"90",
		X"CD",X"3C",X"56",X"DD",X"21",X"E8",X"61",X"21",X"01",X"92",X"06",X"01",X"CD",X"41",X"56",X"DD",
		X"21",X"E9",X"61",X"21",X"C1",X"91",X"06",X"01",X"CD",X"41",X"56",X"C9",X"06",X"03",X"11",X"20",
		X"00",X"DD",X"7E",X"00",X"CD",X"4D",X"56",X"DD",X"23",X"19",X"10",X"F5",X"C9",X"F5",X"E6",X"0F",
		X"77",X"19",X"F1",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"E6",X"0F",X"77",X"C9",X"ED",
		X"52",X"06",X"11",X"CD",X"6A",X"56",X"CD",X"75",X"56",X"C9",X"78",X"77",X"E5",X"7C",X"C6",X"08",
		X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"10",X"31",X"3F",X"43",X"52",X"45",X"44",X"49",X"54",X"3F",
		X"10",X"10",X"10",X"48",X"49",X"47",X"48",X"10",X"53",X"43",X"4F",X"52",X"45",X"10",X"10",X"10",
		X"3F",X"47",X"41",X"4D",X"45",X"10",X"4F",X"56",X"45",X"52",X"10",X"3F",X"10",X"10",X"10",X"10",
		X"10",X"49",X"4E",X"53",X"45",X"52",X"54",X"10",X"43",X"30",X"49",X"4E",X"53",X"10",X"10",X"10",
		X"10",X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"50",X"55",X"53",X"48",X"10",X"53",X"54",X"41",
		X"52",X"54",X"10",X"42",X"55",X"54",X"54",X"4F",X"4E",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",
		X"4F",X"4E",X"45",X"10",X"50",X"4C",X"41",X"59",X"45",X"52",X"10",X"4F",X"4E",X"4C",X"59",X"10",
		X"10",X"3F",X"4F",X"4E",X"45",X"10",X"4F",X"52",X"10",X"54",X"57",X"4F",X"10",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"53",X"3F",X"42",X"4F",X"4E",X"55",X"53",X"3F",X"56",X"41",X"4C",X"41",X"44",
		X"4F",X"4E",X"10",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",X"49",X"4F",X"4E",X"3F",X"10",X"10",
		X"10",X"10",X"10",X"10",X"4D",X"4F",X"56",X"45",X"10",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",
		X"4B",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"54",X"4F",X"10",X"44",X"49",X"53",X"50",
		X"4C",X"41",X"59",X"10",X"59",X"4F",X"55",X"52",X"10",X"4E",X"41",X"4D",X"45",X"10",X"3F",X"53",
		X"43",X"4F",X"52",X"45",X"3F",X"4E",X"41",X"4D",X"45",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"10",X"31",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",X"10",X"32",X"3F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"45",X"4E",X"44",X"10",X"42",X"59",X"10",X"41",X"43",
		X"54",X"49",X"4F",X"4E",X"10",X"42",X"55",X"54",X"54",X"4F",X"4E",X"10",X"10",X"10",X"3F",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"10",X"31",X"39",X"38",X"32",X"3F",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"4A",X"45",X"55",X"10",X"4C",X"45",
		X"10",X"42",X"41",X"47",X"4E",X"41",X"52",X"44",X"3F",X"42",X"52",X"49",X"53",X"53",X"45",X"10",
		X"4A",X"41",X"43",X"51",X"55",X"45",X"53",X"3F",X"37",X"31",X"35",X"33",X"30",X"10",X"43",X"48",
		X"41",X"4C",X"4F",X"4E",X"10",X"53",X"55",X"52",X"10",X"53",X"41",X"4F",X"4E",X"45",X"3F",X"46",
		X"52",X"41",X"4E",X"43",X"45",X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",X"31",X"3F",X"43",
		X"52",X"45",X"44",X"49",X"54",X"3F",X"4D",X"45",X"49",X"4C",X"4C",X"45",X"55",X"52",X"53",X"10",
		X"53",X"43",X"4F",X"52",X"45",X"53",X"3F",X"4A",X"45",X"55",X"10",X"46",X"49",X"4E",X"49",X"10",
		X"10",X"3F",X"49",X"4E",X"54",X"52",X"4F",X"44",X"55",X"49",X"53",X"45",X"5A",X"10",X"56",X"4F",
		X"53",X"10",X"50",X"49",X"45",X"43",X"45",X"53",X"3F",X"41",X"50",X"50",X"55",X"59",X"45",X"5A",
		X"10",X"53",X"55",X"52",X"10",X"4C",X"45",X"10",X"42",X"4F",X"55",X"54",X"4F",X"4E",X"10",X"53",
		X"54",X"41",X"52",X"54",X"3F",X"31",X"10",X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",X"53",X"45",
		X"55",X"4C",X"45",X"4D",X"45",X"4E",X"54",X"3F",X"10",X"10",X"31",X"10",X"4F",X"55",X"10",X"32",
		X"10",X"4A",X"4F",X"55",X"45",X"55",X"52",X"53",X"10",X"10",X"3F",X"42",X"4F",X"4E",X"55",X"53",
		X"3F",X"56",X"41",X"4C",X"41",X"44",X"4F",X"4E",X"10",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",
		X"49",X"4F",X"4E",X"3F",X"55",X"54",X"49",X"4C",X"49",X"53",X"45",X"5A",X"10",X"4C",X"45",X"10",
		X"4D",X"41",X"4E",X"49",X"50",X"55",X"4C",X"41",X"54",X"45",X"55",X"52",X"3F",X"50",X"4F",X"55",
		X"52",X"10",X"49",X"4E",X"53",X"43",X"52",X"49",X"52",X"45",X"10",X"56",X"4F",X"54",X"52",X"45",
		X"10",X"4E",X"4F",X"4D",X"3F",X"53",X"43",X"4F",X"52",X"45",X"3F",X"4E",X"4F",X"4D",X"10",X"3F",
		X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",X"31",X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",
		X"32",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"41",X"43",
		X"54",X"49",X"4F",X"4E",X"10",X"50",X"4F",X"55",X"52",X"10",X"46",X"49",X"4E",X"49",X"52",X"10",
		X"10",X"10",X"10",X"10",X"3F",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"10",X"31",
		X"39",X"38",X"32",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",
		X"80",X"40",X"20",X"10",X"40",X"C4",X"E0",X"40",X"CA",X"D0",X"42",X"E4",X"A0",X"42",X"EA",X"B0",
		X"42",X"EE",X"B0",X"42",X"F0",X"70",X"42",X"F5",X"B0",X"43",X"70",X"B0",X"43",X"78",X"90",X"41",
		X"6F",X"60",X"41",X"74",X"D0",X"42",X"F8",X"70",X"42",X"FA",X"B0",X"42",X"FE",X"D0",X"44",X"87",
		X"E0",X"44",X"8F",X"D0",X"45",X"27",X"A0",X"45",X"2C",X"90",X"45",X"4F",X"80",X"44",X"B3",X"80",
		X"45",X"13",X"40",X"45",X"19",X"60",X"45",X"1B",X"B0",X"45",X"1E",X"D0",X"45",X"AA",X"40",X"46",
		X"CA",X"D0",X"47",X"6A",X"E0",X"47",X"6E",X"90",X"46",X"73",X"E0",X"46",X"78",X"B0",X"46",X"7E",
		X"D0",X"46",X"C4",X"E0",X"48",X"E4",X"E0",X"48",X"87",X"60",X"48",X"8B",X"50",X"48",X"EB",X"E0",
		X"4A",X"27",X"E0",X"4A",X"2B",X"90",X"48",X"F4",X"D0",X"48",X"94",X"60",X"48",X"9B",X"50",X"49",
		X"D1",X"60",X"49",X"D4",X"90",X"49",X"D7",X"E0",X"49",X"DB",X"D0",X"4A",X"E7",X"80",X"4A",X"F0",
		X"80",X"4A",X"F7",X"80",X"4B",X"47",X"40",X"4B",X"53",X"40",X"48",X"E7",X"D0",X"FF",X"FF",X"FF",
		X"40",X"C4",X"80",X"40",X"CA",X"80",X"42",X"E4",X"80",X"42",X"EA",X"80",X"42",X"EE",X"10",X"42",
		X"F0",X"10",X"42",X"F5",X"10",X"43",X"70",X"80",X"43",X"78",X"80",X"41",X"6F",X"40",X"41",X"74",
		X"40",X"42",X"F8",X"20",X"42",X"FA",X"20",X"42",X"FE",X"80",X"FF",X"FF",X"FF",X"44",X"87",X"20",
		X"44",X"8F",X"40",X"45",X"27",X"80",X"45",X"2C",X"10",X"45",X"4F",X"40",X"44",X"B3",X"40",X"45",
		X"13",X"40",X"45",X"19",X"20",X"45",X"1B",X"20",X"45",X"1E",X"40",X"45",X"AA",X"40",X"46",X"CA",
		X"40",X"47",X"6A",X"40",X"47",X"6E",X"10",X"46",X"73",X"20",X"46",X"78",X"20",X"46",X"7E",X"40",
		X"46",X"C4",X"40",X"FF",X"FF",X"FF",X"44",X"87",X"80",X"44",X"8F",X"10",X"45",X"27",X"80",X"45",
		X"2C",X"10",X"45",X"4F",X"80",X"44",X"B3",X"80",X"45",X"13",X"80",X"45",X"19",X"80",X"45",X"1B",
		X"80",X"45",X"1E",X"10",X"45",X"AA",X"80",X"46",X"CA",X"10",X"47",X"6A",X"80",X"47",X"6E",X"10",
		X"46",X"73",X"20",X"46",X"78",X"20",X"46",X"7E",X"80",X"FF",X"FF",X"FF",X"46",X"C4",X"20",X"48",
		X"E4",X"20",X"48",X"87",X"20",X"48",X"8B",X"40",X"48",X"EB",X"20",X"4A",X"27",X"20",X"4A",X"2B",
		X"80",X"48",X"F4",X"80",X"48",X"94",X"20",X"48",X"9B",X"40",X"49",X"D1",X"20",X"49",X"D4",X"80",
		X"49",X"D7",X"20",X"49",X"DB",X"40",X"4A",X"E7",X"80",X"4A",X"F0",X"80",X"4A",X"F7",X"80",X"4B",
		X"47",X"40",X"4B",X"53",X"40",X"FF",X"FF",X"FF",X"58",X"93",X"02",X"A8",X"91",X"01",X"12",X"91",
		X"01",X"98",X"90",X"01",X"2E",X"93",X"01",X"36",X"93",X"01",X"C8",X"91",X"02",X"4C",X"92",X"02",
		X"CA",X"90",X"02",X"CD",X"90",X"02",X"91",X"90",X"02",X"9C",X"90",X"02",X"62",X"90",X"03",X"65",
		X"91",X"03",X"69",X"91",X"03",X"15",X"92",X"03",X"99",X"92",X"03",X"39",X"91",X"03",X"F1",X"F2",
		X"F3",X"F4",X"F5",X"F6",X"F7",X"1F",X"1F",X"1F",X"FF",X"09",X"00",X"1F",X"1F",X"1F",X"FF",X"02",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"20",X"00",X"00",X"03",X"00",X"00",X"00",X"15",
		X"1B",X"00",X"00",X"0C",X"1B",X"00",X"00",X"0C",X"1B",X"00",X"00",X"0C",X"1C",X"00",X"00",X"0C",
		X"1B",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"1F",X"00",X"00",X"16",X"20",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"24",X"19",X"00",X"0C",X"20",X"1A",X"00",X"0C",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"1B",X"00",X"00",X"0C",X"20",X"00",X"00",X"0C",
		X"24",X"00",X"00",X"0C",X"27",X"00",X"00",X"0C",X"24",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"FF",X"1B",X"00",X"00",X"0C",X"20",X"00",X"00",X"0C",X"24",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"1B",X"0F",X"00",X"02",X"18",X"0E",X"00",X"0C",
		X"14",X"0E",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"7F",X"75",X"CE",X"99",
		X"C0",X"8B",X"C4",X"82",X"65",X"96",X"01",X"9E",X"65",X"8B",X"B4",X"8D",X"B0",X"CB",X"3F",X"CB",
		X"3F",X"FE",X"00",X"CA",X"C2",X"55",X"C3",X"B8",X"55",X"20",X"00",X"00",X"02",X"00",X"00",X"00",
		X"08",X"1B",X"00",X"00",X"0F",X"1B",X"00",X"00",X"08",X"1B",X"00",X"00",X"08",X"1C",X"00",X"00",
		X"08",X"00",X"00",X"00",X"08",X"1B",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"1F",X"00",X"00",
		X"20",X"20",X"00",X"00",X"0F",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"FF",X"FF",X"08",X"00",
		X"3A",X"F5",X"61",X"FE",X"00",X"C2",X"68",X"05",X"3A",X"CF",X"61",X"FE",X"00",X"C2",X"68",X"05",
		X"C3",X"5B",X"05",X"26",X"3A",X"F5",X"61",X"FE",X"00",X"C2",X"52",X"06",X"3A",X"CF",X"61",X"FE",
		X"00",X"C2",X"52",X"06",X"C3",X"45",X"06",X"05",X"50",X"50",X"49",X"60",X"46",X"44",X"0C",X"04",
		X"3A",X"59",X"61",X"FE",X"01",X"C8",X"3A",X"5E",X"61",X"FE",X"01",X"C8",X"0A",X"D9",X"FE",X"00",
		X"C3",X"AE",X"23",X"FF",X"58",X"93",X"02",X"A8",X"91",X"01",X"12",X"91",X"01",X"98",X"90",X"01",
		X"DC",X"91",X"01",X"36",X"93",X"01",X"71",X"90",X"01",X"4C",X"92",X"02",X"CA",X"90",X"02",X"C5",
		X"90",X"02",X"91",X"90",X"02",X"9C",X"90",X"02",X"71",X"93",X"03",X"85",X"92",X"03",X"C9",X"91",
		X"03",X"15",X"92",X"03",X"99",X"92",X"03",X"F9",X"90",X"03",X"FF",X"10",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"54",X"60",X"FE",X"00",X"C8",X"CD",X"00",X"55",X"C9",X"C3",X"46",X"5E",X"FE",X"01",X"C8",
		X"DD",X"21",X"44",X"5D",X"FD",X"21",X"80",X"65",X"11",X"04",X"00",X"3A",X"88",X"62",X"FE",X"00",
		X"CC",X"2A",X"5D",X"3A",X"88",X"62",X"FE",X"00",X"28",X"05",X"DD",X"19",X"3D",X"18",X"F7",X"DD",
		X"7E",X"03",X"FE",X"FF",X"28",X"3C",X"FE",X"FE",X"CA",X"1C",X"5D",X"47",X"3A",X"26",X"60",X"E6",
		X"07",X"B0",X"32",X"26",X"60",X"FD",X"7E",X"02",X"DD",X"BE",X"00",X"C0",X"FD",X"7E",X"03",X"DD",
		X"BE",X"01",X"C0",X"3A",X"0D",X"60",X"DD",X"BE",X"02",X"C0",X"3A",X"88",X"62",X"3C",X"32",X"88",
		X"62",X"3A",X"26",X"60",X"E6",X"80",X"FE",X"80",X"C8",X"3A",X"26",X"60",X"E6",X"07",X"32",X"26",
		X"60",X"C9",X"3E",X"10",X"32",X"97",X"65",X"32",X"9B",X"65",X"3E",X"D0",X"32",X"96",X"65",X"3E",
		X"E0",X"C3",X"38",X"5E",X"3A",X"87",X"65",X"FE",X"11",X"C0",X"18",X"CE",X"3A",X"8A",X"65",X"FE",
		X"7F",X"C0",X"3A",X"19",X"60",X"FE",X"01",X"C0",X"18",X"C0",X"21",X"C2",X"91",X"22",X"C4",X"61",
		X"22",X"FA",X"61",X"3E",X"01",X"32",X"C6",X"61",X"32",X"FC",X"61",X"3E",X"03",X"32",X"99",X"60",
		X"32",X"9A",X"60",X"C9",X"3C",X"E0",X"01",X"10",X"3C",X"70",X"01",X"20",X"28",X"70",X"01",X"08",
		X"28",X"70",X"01",X"80",X"28",X"70",X"01",X"00",X"28",X"70",X"01",X"00",X"28",X"70",X"01",X"00",
		X"39",X"70",X"01",X"10",X"3C",X"11",X"01",X"20",X"85",X"10",X"01",X"10",X"85",X"10",X"01",X"80",
		X"85",X"10",X"01",X"00",X"85",X"10",X"01",X"00",X"85",X"10",X"01",X"00",X"56",X"10",X"01",X"08",
		X"7D",X"10",X"01",X"10",X"7D",X"10",X"01",X"80",X"7D",X"10",X"01",X"00",X"7D",X"10",X"01",X"00",
		X"7D",X"10",X"01",X"00",X"6C",X"10",X"02",X"10",X"6C",X"10",X"02",X"80",X"6C",X"10",X"02",X"00",
		X"6C",X"10",X"02",X"00",X"6C",X"10",X"02",X"00",X"8C",X"10",X"02",X"10",X"8C",X"10",X"02",X"FF",
		X"98",X"10",X"02",X"10",X"98",X"88",X"02",X"00",X"38",X"88",X"02",X"08",X"38",X"88",X"02",X"80",
		X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",
		X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",
		X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",
		X"5B",X"88",X"02",X"10",X"5C",X"C0",X"02",X"40",X"40",X"C0",X"02",X"08",X"44",X"C0",X"02",X"10",
		X"40",X"C0",X"02",X"08",X"44",X"C0",X"02",X"10",X"40",X"C0",X"02",X"08",X"59",X"C0",X"02",X"10",
		X"5C",X"E0",X"02",X"40",X"7D",X"E0",X"02",X"10",X"7D",X"E0",X"02",X"80",X"7D",X"E0",X"02",X"FE",
		X"7D",X"E0",X"02",X"80",X"B9",X"E0",X"02",X"00",X"B4",X"C8",X"02",X"20",X"B8",X"C8",X"02",X"10",
		X"FF",X"FF",X"FF",X"10",X"60",X"FF",X"FF",X"FF",X"32",X"9A",X"65",X"3E",X"03",X"32",X"99",X"60",
		X"32",X"9A",X"60",X"C3",X"14",X"5D",X"3A",X"54",X"60",X"FE",X"01",X"C8",X"3A",X"26",X"60",X"E6",
		X"07",X"32",X"26",X"60",X"C3",X"A0",X"5C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"0A",X"32",X"7D",X"62",X"0E",X"01",X"C9",X"FF",X"32",X"ED",X"61",X"3E",X"0A",X"32",X"7D",
		X"62",X"C3",X"C9",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"18",X"0C",X"1C",X"5C",X"F8",
		X"60",X"74",X"7D",X"79",X"3E",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"EC",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"1C",X"1F",X"1F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"60",X"F8",X"F8",X"F8",X"F0",
		X"7F",X"7F",X"7F",X"1B",X"03",X"01",X"00",X"00",X"F0",X"FC",X"FC",X"FC",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"74",X"00",X"00",X"00",X"18",X"0C",X"5C",X"DC",X"F8",
		X"7D",X"79",X"3E",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"EC",X"C0",X"80",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"3F",X"3F",X"3F",X"07",X"0F",X"1F",X"07",X"0F",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"03",X"0F",
		X"04",X"04",X"00",X"20",X"70",X"21",X"00",X"80",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"0F",X"8F",
		X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"EF",X"FF",X"0F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"00",X"00",X"18",X"3C",X"3C",X"3C",X"3F",
		X"07",X"07",X"06",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"7E",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"7C",X"FC",
		X"3F",X"3F",X"79",X"3E",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"60",X"75",X"7D",X"79",X"3E",X"00",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"07",X"07",X"07",X"0F",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"3F",X"07",X"47",X"C3",X"EB",X"FB",X"F2",X"7C",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1D",X"00",X"00",X"00",X"70",X"70",X"E0",X"E0",X"EC",
		X"0F",X"07",X"43",X"C1",X"E9",X"FB",X"F6",X"7C",X"F8",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C1",X"00",X"00",X"00",X"00",X"38",X"78",X"F8",X"F0",
		X"E9",X"FB",X"F3",X"7D",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"F8",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"3A",X"00",X"00",X"00",X"00",X"08",X"1C",X"3C",X"7C",
		X"3E",X"3C",X"1F",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"78",X"7C",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"0C",X"1C",X"DC",X"F8",
		X"74",X"7D",X"79",X"3E",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"4C",X"5C",
		X"74",X"7D",X"79",X"3E",X"00",X"00",X"00",X"00",X"D8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"3F",X"3F",X"3F",X"07",X"0F",X"1F",X"07",X"07",
		X"02",X"20",X"70",X"20",X"00",X"04",X"0E",X"04",X"07",X"03",X"00",X"06",X"02",X"07",X"7F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"3F",X"3F",X"3F",X"07",X"07",X"0F",X"03",X"0F",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"03",X"00",X"06",X"02",X"07",X"7F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"07",X"0F",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"06",X"02",X"07",X"7F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"3F",X"3F",X"07",X"0F",X"8F",X"8F",X"8F",
		X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"CF",X"FF",X"3F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"0C",X"00",X"00",X"00",X"18",X"1C",X"3C",X"3C",X"3F",
		X"07",X"07",X"0F",X"07",X"01",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"FF",X"FE",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"7C",X"FC",
		X"3F",X"3F",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"1F",X"1F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"F0",
		X"7F",X"7F",X"7F",X"1B",X"03",X"01",X"00",X"00",X"F0",X"FC",X"FC",X"FC",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"00",X"00",X"10",X"18",X"1C",X"0C",X"5C",X"D8",
		X"60",X"74",X"70",X"71",X"3E",X"08",X"00",X"00",X"FC",X"FC",X"FC",X"EC",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"74",X"00",X"00",X"10",X"18",X"1C",X"4C",X"DC",X"D8",
		X"7D",X"71",X"3E",X"08",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"E0",X"C0",X"80",X"00",X"00",
		X"08",X"04",X"02",X"01",X"20",X"20",X"20",X"60",X"00",X"00",X"00",X"00",X"08",X"3C",X"FC",X"FC",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"80",X"80",X"5C",X"FC",X"FC",
		X"60",X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"F8",X"F8",X"FC",X"FC",X"F8",X"68",X"00",X"00",
		X"08",X"04",X"02",X"01",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"08",X"1C",X"7C",X"FC",
		X"60",X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"F8",X"F8",X"FC",X"FC",X"F8",X"68",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"20",X"20",X"20",X"00",X"28",X"1C",X"FC",X"FC",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"3A",X"10",X"10",X"10",X"00",X"18",X"1C",X"3C",X"7C",
		X"3E",X"38",X"1F",X"07",X"01",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"7C",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"80",X"80",X"80",X"00",X"9C",X"3C",X"7C",X"F8",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"F8",X"FC",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"40",X"40",X"40",X"00",X"4C",X"1C",X"DC",X"F8",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"00",X"00",X"00",X"10",X"18",X"3C",X"4C",X"DC",
		X"74",X"70",X"71",X"3E",X"0E",X"02",X"00",X"00",X"D8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"00",X"09",X"25",X"D4",X"B5",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"02",X"03",X"01",X"07",X"0F",X"0D",X"08",X"00",X"1C",X"7E",X"A3",X"FF",X"AB",X"FF",X"AB",X"8B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"08",X"08",X"0E",X"0F",X"0E",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0E",X"0F",X"0E",X"08",X"08",X"1C",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1C",X"1E",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"9F",X"8F",X"8F",X"87",X"83",X"81",X"80",
		X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"BF",
		X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"87",X"87",X"87",X"87",X"83",X"83",X"83",X"83",
		X"9F",X"9F",X"8F",X"8F",X"8F",X"8F",X"8F",X"87",X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",
		X"9F",X"9F",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"8F",X"8F",X"8F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"81",X"83",X"83",X"87",X"87",X"87",X"8F",X"8F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"9F",X"8F",X"87",X"87",X"83",X"81",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"87",X"83",X"83",X"81",X"81",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"8F",X"8F",X"8F",X"8F",X"87",X"87",X"87",X"87",X"8F",X"8F",X"8F",X"8F",X"9F",X"9F",X"9F",
		X"80",X"80",X"81",X"81",X"83",X"83",X"87",X"87",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"B8",X"B0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"BF",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"0C",X"10",X"30",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"26",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"64",X"74",X"7C",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"3A",X"18",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"64",X"74",X"7C",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"3A",X"09",X"08",X"08",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"01",X"01",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"A0",X"B8",X"B4",X"EA",X"AE",X"9A",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"10",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"10",X"30",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"70",X"70",X"70",X"70",X"70",X"70",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"03",X"06",X"0C",X"18",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F8",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"3C",X"7E",X"FF",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"FF",X"7E",X"3C",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"01",X"03",X"07",X"1F",X"1F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"0E",X"1E",X"1E",
		X"1E",X"1E",X"1E",X"10",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",
		X"00",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"00",X"10",X"18",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"47",X"57",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"18",X"00",X"00",X"00",
		X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"18",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"04",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"18",X"00",X"00",X"00",X"00",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"18",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"18",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"04",X"00",X"00",X"10",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"02",X"00",X"00",X"00",X"00",X"08",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"06",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"02",X"00",X"00",X"00",X"00",X"08",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"06",X"06",X"06",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"71",X"89",X"89",X"89",X"89",X"89",X"67",X"00",X"6E",X"91",X"91",X"91",X"91",X"91",X"6E",X"00",
		X"7E",X"91",X"91",X"91",X"91",X"91",X"61",X"00",X"FF",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"C3",X"A5",X"A5",X"A5",X"BD",X"C3",X"7E",X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",
		X"00",X"7F",X"02",X"04",X"08",X"10",X"20",X"7F",X"00",X"06",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",
		X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"8F",X"2F",X"EF",X"EF",X"EF",X"EF",X"8F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E3",
		X"8F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"37",X"77",X"77",X"37",X"87",X"E7",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"F8",X"F3",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F3",X"F8",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"2F",X"0F",X"7F",X"7F",
		X"3F",X"8F",X"E7",X"F7",X"F7",X"F7",X"F7",X"F7",X"0F",X"EF",X"EF",X"EF",X"CF",X"DF",X"DF",X"9F",
		X"87",X"BF",X"BF",X"BF",X"9F",X"DF",X"DF",X"CF",X"BF",X"BF",X"3F",X"7F",X"7F",X"7F",X"0F",X"EF",
		X"EF",X"EF",X"E7",X"F7",X"F7",X"F7",X"87",X"BF",X"EF",X"0F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"1F",X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"8F",X"1F",X"7F",X"FF",
		X"BF",X"87",X"F7",X"77",X"17",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"C7",X"F1",X"FC",X"FE",X"FE",
		X"FC",X"F1",X"C7",X"1F",X"7F",X"FF",X"FC",X"F9",X"C7",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F1",X"F4",X"F7",X"F7",X"F7",X"F7",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",X"F7",X"F7",X"F7",X"F7",X"F4",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"80",X"41",X"AA",X"00",X"00",X"00",X"02",X"15",X"2A",X"55",X"AA",
		X"00",X"00",X"00",X"80",X"40",X"A8",X"55",X"AA",X"01",X"02",X"15",X"AA",X"55",X"AA",X"55",X"AA",
		X"40",X"80",X"50",X"A8",X"55",X"AA",X"55",X"AA",X"15",X"2A",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"50",X"A8",X"54",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"07",
		X"F0",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"03",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"FC",X"FC",X"FC",X"FC",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"00",X"01",X"01",X"01",X"00",X"00",X"10",X"10",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"78",X"38",X"00",X"00",X"10",X"10",X"1F",X"3F",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"1C",X"1E",X"1F",X"1F",X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"01",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7E",X"7C",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"7F",X"7F",X"7F",X"7F",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"01",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",
		X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"10",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"C0",X"FF",X"FF",X"FE",X"FE",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"00",X"00",X"10",X"10",
		X"80",X"80",X"80",X"80",X"00",X"00",X"10",X"10",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"0F",X"0F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",
		X"01",X"03",X"03",X"07",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"FE",X"FE",X"FF",X"FF",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"FE",X"FE",X"FF",X"FF",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"7F",X"3F",X"1F",X"0F",X"07",X"07",X"03",X"01",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"FF",X"7F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"00",X"01",X"03",X"03",X"07",X"0F",X"0F",X"1F",
		X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1E",X"1C",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"3F",X"3F",X"3F",X"7F",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",
		X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"60",X"20",X"00",X"00",X"10",X"10",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"0E",X"0C",X"00",X"00",X"10",X"10",
		X"00",X"00",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",
		X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FC",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",
		X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FE",X"FE",X"FE",X"00",X"00",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"F0",X"F8",X"F8",X"FC",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"00",X"00",X"00",X"09",X"3B",X"2B",X"2B",X"A8",
		X"7F",X"6B",X"62",X"46",X"00",X"07",X"06",X"00",X"A9",X"AB",X"AB",X"AB",X"80",X"80",X"00",X"00",
		X"00",X"00",X"C8",X"EA",X"02",X"42",X"62",X"60",X"00",X"00",X"00",X"20",X"A8",X"A8",X"A8",X"A0",
		X"60",X"62",X"42",X"02",X"02",X"00",X"00",X"00",X"A1",X"AB",X"AB",X"AA",X"A0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"6B",X"00",X"00",X"00",X"09",X"3B",X"2B",X"AB",X"A8",
		X"62",X"46",X"01",X"07",X"07",X"03",X"00",X"00",X"A9",X"AB",X"AB",X"AB",X"80",X"80",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"D7",X"D0",X"D7",X"80",X"0F",X"20",X"3F",X"00",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"00",X"3F",X"D0",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"A0",X"AE",X"12",X"0A",X"0A",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"1F",X"00",X"00",X"00",X"11",X"17",X"97",X"07",X"05",
		X"1D",X"1D",X"01",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"D5",X"54",X"54",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"FF",X"00",X"00",X"00",X"00",X"09",X"2B",X"2B",X"AB",
		X"EA",X"EA",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A9",X"AB",X"AB",X"2B",X"00",X"00",X"00",
		X"00",X"03",X"01",X"00",X"01",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"0C",X"36",X"7F",X"6B",X"62",X"46",X"00",X"00",X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"00",X"07",X"00",X"0F",X"80",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"E8",X"1F",X"68",X"FF",X"D4",X"C7",X"8C",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"70",X"75",X"00",X"F0",X"70",X"00",X"70",X"40",X"40",X"41",
		X"05",X"1D",X"6D",X"FF",X"D5",X"C5",X"8C",X"00",X"57",X"57",X"56",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"6C",X"FE",X"00",X"00",X"78",X"B8",X"90",X"D0",X"50",X"50",
		X"D7",X"C5",X"8D",X"01",X"00",X"00",X"01",X"00",X"50",X"50",X"50",X"50",X"50",X"90",X"B8",X"3C",
		X"00",X"00",X"00",X"00",X"06",X"1B",X"3F",X"35",X"00",X"00",X"00",X"30",X"20",X"35",X"97",X"D7",
		X"31",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"53",X"50",X"50",X"54",X"54",X"54",X"DC",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"00",X"00",X"3C",X"DC",X"88",X"88",X"88",X"A8",
		X"6B",X"62",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A8",X"A8",X"A9",X"2F",X"2F",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"00",X"00",X"00",X"00",X"09",X"2B",X"3B",X"AB",
		X"6B",X"62",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A9",X"AB",X"AB",X"2B",X"00",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"C0",X"C0",X"C0",X"80",X"00",X"3F",X"3F",X"0F",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"C0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"0F",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"10",X"38",X"5C",
		X"02",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"7C",X"FC",X"FE",X"FF",X"FF",X"3F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"13",X"00",X"00",X"00",X"01",X"03",X"23",X"F3",X"F0",
		X"1F",X"1F",X"07",X"07",X"01",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"9F",X"00",X"00",X"00",X"00",X"01",X"23",X"63",X"E3",
		X"FF",X"FF",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E1",X"E3",X"E3",X"63",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"FF",X"1F",X"3D",X"1C",X"1E",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"00",
		X"1E",X"1C",X"3D",X"1B",X"03",X"01",X"00",X"00",X"01",X"83",X"83",X"82",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"16",X"00",X"00",X"10",X"11",X"13",X"33",X"33",X"20",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0F",X"06",X"00",X"E1",X"F3",X"F3",X"E3",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"1F",X"00",X"00",X"10",X"11",X"13",X"73",X"F3",X"E0",
		X"10",X"3F",X"3E",X"0E",X"07",X"03",X"00",X"00",X"E1",X"F3",X"F3",X"E3",X"C0",X"80",X"00",X"00",
		X"08",X"04",X"02",X"01",X"04",X"0C",X"16",X"1F",X"00",X"00",X"00",X"80",X"C0",X"61",X"E3",X"E3",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C3",X"C0",X"E0",X"E1",X"67",X"07",X"06",X"00",
		X"00",X"00",X"00",X"1F",X"01",X"04",X"0C",X"16",X"00",X"00",X"00",X"80",X"80",X"C1",X"E3",X"E3",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"E3",X"C0",X"C0",X"E1",X"E7",X"67",X"06",X"00",
		X"08",X"04",X"02",X"01",X"00",X"04",X"0C",X"16",X"00",X"00",X"00",X"80",X"C0",X"41",X"63",X"E3",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"E3",X"C0",X"C0",X"E1",X"E7",X"67",X"06",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"20",X"20",X"20",X"60",X"60",X"41",X"E3",X"E3",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C3",X"C0",X"E0",X"E1",X"67",X"07",X"06",X"00",
		X"00",X"00",X"00",X"02",X"06",X"0B",X"0F",X"0F",X"10",X"10",X"10",X"30",X"30",X"21",X"B3",X"F3",
		X"0F",X"1F",X"1F",X"07",X"01",X"00",X"00",X"00",X"F3",X"E0",X"E0",X"60",X"60",X"40",X"DC",X"DE",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"00",X"80",X"BC",X"DC",X"C0",X"60",X"60",X"E0",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E0",X"E0",X"60",X"40",X"DC",X"DE",X"DE",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"40",X"40",X"7C",X"DC",X"C0",X"80",X"C0",X"C0",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C0",X"C0",X"E0",X"E1",X"67",X"27",X"66",X"60",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"00",X"00",X"00",X"10",X"11",X"13",X"33",X"33",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E1",X"F3",X"F3",X"63",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"00",X"00",X"0E",X"8C",X"CC",X"EA",X"00",X"00",X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",X"FE",X"54",X"FE",X"54",X"74",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"C8",X"E8",X"F2",X"F3",X"F2",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F2",X"F3",X"F2",X"E8",X"C8",X"9C",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"01",X"01",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"07",X"02",X"02",X"02",X"02",X"02",X"02",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"A0",X"A0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"BE",X"BF",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"A0",X"80",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"A0",X"A0",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",X"80",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"BF",X"BF",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"BC",X"BC",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B8",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"A0",X"A0",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"A0",X"A0",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"B0",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"BC",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"9F",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"BF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"B8",X"B8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"A0",X"A0",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"B8",X"B8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",
		X"8F",X"9F",X"BF",X"BF",X"FF",X"FF",X"BF",X"BF",X"80",X"81",X"81",X"83",X"83",X"87",X"87",X"8F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"81",X"81",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"1F",X"0E",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"14",X"0C",X"0C",X"0A",X"18",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0F",X"0F",X"0E",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0C",X"0C",X"0A",X"09",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"D8",X"5C",X"76",X"74",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"75",
		X"7A",X"35",X"3A",X"15",X"1A",X"05",X"0A",X"05",X"1A",X"15",X"1A",X"15",X"0A",X"05",X"0A",X"05",
		X"FA",X"F5",X"7A",X"75",X"7A",X"35",X"3A",X"35",X"FA",X"F5",X"FA",X"75",X"7A",X"35",X"3A",X"15",
		X"EA",X"E5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"8A",X"85",X"8A",X"85",X"8A",X"85",
		X"8A",X"85",X"8A",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"EA",X"E5",X"EA",X"E5",X"EA",X"E5",
		X"7A",X"75",X"7A",X"75",X"FA",X"F5",X"FA",X"F5",X"1A",X"15",X"3A",X"35",X"3A",X"35",X"7A",X"75",
		X"7A",X"75",X"7A",X"75",X"3A",X"35",X"3A",X"35",X"3A",X"35",X"3A",X"35",X"7A",X"75",X"7A",X"75",
		X"EA",X"C5",X"CA",X"85",X"8A",X"05",X"0A",X"05",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"E5",
		X"0A",X"85",X"CA",X"E5",X"FA",X"F5",X"FA",X"F5",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",
		X"FA",X"F5",X"FA",X"E5",X"EA",X"E5",X"CA",X"C5",X"CA",X"C5",X"8A",X"85",X"8A",X"85",X"8A",X"85",
		X"8A",X"85",X"8A",X"85",X"8A",X"85",X"8A",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"EA",X"E5",
		X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"1A",X"15",X"1A",X"15",X"3A",X"75",X"7A",X"75",
		X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"FF",X"04",X"08",X"10",X"20",X"40",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"40",X"A0",X"50",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"A0",X"50",X"A0",X"40",X"A0",X"50",X"A0",X"50",X"AF",X"5F",X"AF",X"5F",X"AF",X"FF",X"FF",X"FF",
		X"04",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1A",
		X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"20",X"20",X"3E",X"20",X"20",
		X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"02",X"02",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"2E",X"2A",X"2A",X"2A",X"3A",
		X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",X"2A",X"2A",
		X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"20",X"3E",X"20",X"20",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",
		X"00",X"3E",X"10",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"20",X"1E",X"24",X"24",X"24",X"1E",X"00",X"20",X"28",X"28",X"28",X"3E",X"00",X"20",
		X"28",X"28",X"28",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",
		X"3E",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",
		X"02",X"04",X"38",X"00",X"1C",X"22",X"22",X"22",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",X"3E",X"00",
		X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",X"02",X"04",
		X"38",X"00",X"1E",X"24",X"24",X"24",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",
		X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",
		X"20",X"20",X"3E",X"20",X"20",X"00",X"3E",X"00",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",
		X"22",X"22",X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"20",X"20",X"3E",
		X"20",X"20",X"00",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"38",X"04",X"02",X"3C",X"02",
		X"08",X"08",X"08",X"08",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"E0",X"30",X"18",X"08",X"08",X"08",X"08",X"08",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F8",X"E4",X"E2",X"E2",X"E2",X"E3",X"E3",X"FE",X"E0",X"0E",X"31",X"61",X"E1",
		X"E1",X"E1",X"E1",X"EE",X"F0",X"E0",X"FE",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"FC",X"00",
		X"F8",X"E6",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"EE",X"F0",X"E0",X"E0",X"F0",X"E8",X"E4",
		X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"72",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"07",X"04",X"02",X"01",X"02",X"04",X"07",
		X"00",X"04",X"04",X"07",X"04",X"04",X"E0",X"FC",X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",
		X"FC",X"E0",X"80",X"00",X"FC",X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E6",X"F8",X"00",X"F8",
		X"E6",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"EC",X"F0",X"E0",X"E0",X"E0",X"F8",X"E4",
		X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"7B",X"06",X"E0",X"FC",X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"E2",X"FE",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"EC",X"E2",X"E3",X"E3",X"E3",X"E3",
		X"E3",X"E3",X"E6",X"E8",X"00",X"E0",X"E8",X"E4",X"E2",X"E2",X"E2",X"E3",X"E3",X"63",X"63",X"63",
		X"63",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"E2",X"E2",X"EC",X"F0",X"00",X"F8",X"E6",X"E3",X"E3",
		X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"EC",X"F0",X"E0",X"E0",X"E0",X"E8",X"E4",X"E2",X"E2",X"E3",
		X"E3",X"E3",X"E3",X"7B",X"06",X"E0",X"E8",X"E4",X"E2",X"E3",X"E3",X"E3",X"E3",X"23",X"23",X"23",
		X"23",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"E2",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"11",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"FF",X"00",X"00",
		X"07",X"19",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"FD",X"F3",X"E1",X"F1",X"F9",X"F7",X"F1",X"F1",
		X"F1",X"F1",X"71",X"19",X"07",X"01",X"00",X"00",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"71",X"11",X"11",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"FF",X"00",X"07",X"C9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"C9",X"86",
		X"80",X"C0",X"E1",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"31",X"0E",X"00",X"07",X"19",X"71",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"FD",X"F3",X"E1",X"F1",X"F9",X"F7",X"F1",X"F1",X"F1",X"F1",X"71",
		X"19",X"07",X"01",X"00",X"00",X"01",X"03",X"05",X"05",X"09",X"09",X"C9",X"F1",X"F1",X"F1",X"91",
		X"91",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"07",
		X"00",X"00",X"03",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"06",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",
		X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"06",X"01",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"04",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"02",X"01",X"00",X"01",X"02",X"02",X"04",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"04",X"06",X"01",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"0F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"07",X"07",X"07",X"07",X"87",X"E7",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"20",X"00",X"00",X"00",
		X"3F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"07",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"3F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"3F",X"07",X"07",X"07",X"07",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"07",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"12",X"01",X"00",X"22",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"50",X"00",X"00",X"00",X"00",X"02",X"15",X"2A",X"55",
		X"00",X"00",X"00",X"00",X"80",X"40",X"A8",X"55",X"00",X"01",X"02",X"15",X"AA",X"55",X"AA",X"55",
		X"80",X"40",X"80",X"50",X"A8",X"55",X"AA",X"55",X"0A",X"15",X"2A",X"55",X"AA",X"55",X"AA",X"55",
		X"0A",X"50",X"A8",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",
		X"0F",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"03",X"01",X"01",X"01",X"00",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"01",X"01",X"00",X"00",X"03",X"03",X"03",X"03",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"10",X"10",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"00",X"00",X"10",X"10",X"E0",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"07",X"07",X"06",X"04",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"01",X"01",X"00",X"00",X"7F",X"3F",X"1F",X"1F",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"03",X"03",X"03",X"03",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",
		X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"01",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"03",X"03",X"03",X"01",X"01",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"10",X"10",
		X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"10",X"10",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",
		X"3F",X"3F",X"7F",X"3F",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"F0",X"F0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"FE",X"FC",X"7C",X"38",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"10",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"FC",X"FE",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",
		X"03",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",
		X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"0F",
		X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"FF",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"E0",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"C0",X"C0",X"C0",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"07",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"1F",X"1F",X"00",X"00",X"10",X"10",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",
		X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",
		X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"00",X"00",X"10",X"10",
		X"00",X"00",X"07",X"03",X"01",X"01",X"00",X"00",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"03",
		X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"01",X"01",X"01",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"0C",X"06",X"07",X"03",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		if we = '1' then
			rom_data(to_integer(unsigned(addr))) <= din;
			dout <= din;
		else
			dout <= rom_data(to_integer(unsigned(addr)));
		end if;
	end if;
end process;
end architecture;
