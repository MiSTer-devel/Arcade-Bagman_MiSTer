library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bagman_speech1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bagman_speech1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"E5",X"84",X"FF",X"AC",X"84",X"85",X"85",X"84",X"84",X"84",X"FF",X"FC",X"A5",X"E7",X"B5",
		X"E5",X"A4",X"9F",X"8D",X"FC",X"C5",X"85",X"9C",X"FD",X"E4",X"97",X"ED",X"9F",X"C4",X"A5",X"AF",
		X"D5",X"84",X"84",X"85",X"84",X"84",X"85",X"FE",X"ED",X"B6",X"E5",X"BD",X"A4",X"C5",X"CF",X"F7",
		X"9E",X"C4",X"D5",X"8D",X"8D",X"E4",X"BD",X"87",X"CD",X"C4",X"A4",X"86",X"BD",X"84",X"85",X"84",
		X"84",X"85",X"85",X"FE",X"E4",X"BE",X"D5",X"9C",X"85",X"C7",X"F5",X"EF",X"DD",X"C4",X"8C",X"D4",
		X"95",X"E5",X"BC",X"86",X"D6",X"85",X"E5",X"C7",X"DC",X"85",X"85",X"85",X"84",X"84",X"85",X"FE",
		X"E4",X"9D",X"BC",X"FF",X"84",X"C5",X"FF",X"D6",X"DF",X"C5",X"85",X"DC",X"FC",X"E5",X"8C",X"B7",
		X"AD",X"84",X"E5",X"C7",X"DE",X"84",X"84",X"85",X"84",X"85",X"85",X"FF",X"E5",X"BE",X"9F",X"9D",
		X"84",X"D7",X"EF",X"CC",X"FE",X"D4",X"85",X"8D",X"CD",X"E4",X"95",X"BD",X"A7",X"84",X"D4",X"E7",
		X"BE",X"84",X"85",X"84",X"85",X"84",X"85",X"FF",X"84",X"CF",X"FF",X"FD",X"84",X"CE",X"D7",X"D7",
		X"AD",X"DC",X"84",X"C5",X"B5",X"B4",X"DC",X"EC",X"97",X"84",X"D5",X"EF",X"BF",X"85",X"84",X"85",
		X"85",X"84",X"85",X"FF",X"84",X"D7",X"EC",X"9F",X"85",X"C6",X"DE",X"CF",X"A7",X"DD",X"84",X"E4",
		X"8D",X"BC",X"FC",X"C5",X"CE",X"95",X"C4",X"FF",X"8F",X"84",X"85",X"85",X"85",X"84",X"84",X"FF",
		X"95",X"CF",X"E4",X"8E",X"85",X"D7",X"CE",X"94",X"B4",X"CD",X"94",X"A5",X"87",X"BD",X"CD",X"C7",
		X"A4",X"F4",X"EE",X"ED",X"EC",X"85",X"85",X"84",X"85",X"85",X"84",X"FE",X"BD",X"E7",X"C4",X"94",
		X"84",X"FF",X"F6",X"EC",X"FD",X"E4",X"FD",X"E4",X"F5",X"ED",X"F4",X"F7",X"E7",X"F5",X"FC",X"F6",
		X"FF",X"E4",X"E5",X"E4",X"E4",X"E5",X"E5",X"EE",X"EC",X"F6",X"F7",X"FC",X"E7",X"FD",X"EF",X"E7",
		X"FE",X"F5",X"FD",X"F5",X"FD",X"F5",X"FC",X"FE",X"F6",X"FD",X"FD",X"FE",X"FE",X"F5",X"F5",X"F4",
		X"F4",X"FC",X"FD",X"FE",X"FC",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FC",X"FD",X"FD",X"FD",X"FC",
		X"FC",X"FD",X"FC",X"FF",X"FC",X"FC",X"FF",X"FD",X"FE",X"FC",X"FC",X"FD",X"FC",X"FD",X"FD",X"FF",
		X"FD",X"FE",X"FF",X"FD",X"FF",X"FD",X"FE",X"FD",X"FF",X"FC",X"FD",X"FD",X"FC",X"FC",X"FD",X"FF",
		X"FC",X"FC",X"FE",X"FD",X"FC",X"FC",X"FD",X"FC",X"FD",X"FC",X"FD",X"FF",X"FC",X"FF",X"FF",X"FD",
		X"FE",X"FC",X"FF",X"FD",X"FE",X"FD",X"FC",X"FD",X"FD",X"FC",X"FC",X"FE",X"FF",X"FC",X"FD",X"FF",
		X"FF",X"FD",X"FD",X"FC",X"FC",X"FD",X"FD",X"FE",X"FD",X"FE",X"FE",X"FF",X"FF",X"FE",X"FC",X"FD",
		X"FF",X"FC",X"FC",X"FC",X"FF",X"FC",X"FC",X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",X"FC",X"FD",X"FD",
		X"FD",X"FC",X"FC",X"FF",X"FD",X"FE",X"FF",X"FC",X"FF",X"FD",X"FC",X"FC",X"FE",X"FD",X"FC",X"FD",
		X"FD",X"FD",X"FD",X"FF",X"FC",X"FC",X"FC",X"FF",X"FE",X"FD",X"FD",X"FC",X"FD",X"FD",X"FC",X"FE",
		X"FD",X"FF",X"FE",X"FC",X"FE",X"FF",X"FC",X"FC",X"FF",X"FD",X"FC",X"FC",X"FF",X"FD",X"FC",X"FF",
		X"FD",X"FD",X"FC",X"FE",X"FD",X"FC",X"FC",X"FC",X"FC",X"FD",X"FD",X"FE",X"FC",X"FE",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FD",X"FC",X"FD",X"FF",X"FE",X"FD",X"FE",X"FD",
		X"FC",X"FD",X"FD",X"FC",X"FC",X"FC",X"FD",X"FE",X"FC",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FC",
		X"FF",X"FD",X"FD",X"FC",X"FE",X"FD",X"FC",X"FE",X"FC",X"FC",X"FF",X"FD",X"FC",X"FC",X"FC",X"FD",
		X"FC",X"FD",X"FD",X"FF",X"FD",X"FF",X"FE",X"FC",X"FF",X"FF",X"FE",X"FD",X"FE",X"FC",X"FD",X"FD",
		X"FC",X"FC",X"FD",X"FF",X"FC",X"FC",X"FC",X"FF",X"FE",X"FC",X"FD",X"FD",X"FC",X"FC",X"FD",X"FF",
		X"FC",X"FF",X"FF",X"FD",X"FE",X"FE",X"FD",X"FC",X"FD",X"FD",X"FC",X"FD",X"FD",X"FC",X"FC",X"FE",
		X"FD",X"FC",X"FD",X"FF",X"FF",X"FD",X"FD",X"FC",X"FC",X"FC",X"FD",X"FE",X"FD",X"FE",X"FC",X"FD",
		X"FF",X"FC",X"FC",X"FD",X"FF",X"FC",X"FC",X"FC",X"FD",X"FC",X"FC",X"FF",X"FD",X"FC",X"FE",X"FD",
		X"FD",X"FC",X"FD",X"FD",X"FD",X"FC",X"FC",X"FF",X"FC",X"FF",X"FD",X"FE",X"FF",X"FF",X"FC",X"FE",
		X"FC",X"FD",X"FC",X"FF",X"FF",X"FC",X"FF",X"FD",X"FE",X"FC",X"FC",X"FF",X"FE",X"FD",X"FD",X"FC",
		X"FD",X"FD",X"FC",X"FE",X"FD",X"FD",X"FC",X"FE",X"FC",X"FF",X"FE",X"FC",X"FD",X"FC",X"FD",X"FC",
		X"FD",X"FD",X"FC",X"FF",X"FF",X"FD",X"FE",X"FD",X"FD",X"FC",X"FC",X"FC",X"FC",X"FD",X"FD",X"FE",
		X"FC",X"FE",X"FD",X"FC",X"FF",X"FD",X"FC",X"FD",X"FD",X"FC",X"FC",X"FD",X"FD",X"FC",X"FF",X"FD",
		X"FE",X"FD",X"FF",X"FC",X"FC",X"FD",X"FD",X"FD",X"FC",X"FC",X"FD",X"FF",X"FC",X"FF",X"FC",X"FC",
		X"FE",X"FD",X"FF",X"FC",X"FD",X"FC",X"FD",X"FC",X"FF",X"FD",X"FE",X"FC",X"FC",X"FC",X"FF",X"FD",
		X"FC",X"FC",X"FC",X"FD",X"FC",X"FD",X"FC",X"FF",X"FD",X"FE",X"FD",X"FD",X"FE",X"FF",X"FF",X"FE",
		X"FC",X"FC",X"FD",X"FD",X"FF",X"FC",X"FD",X"FF",X"FF",X"FC",X"FE",X"FD",X"FD",X"FC",X"FD",X"FC",
		X"FD",X"FC",X"FD",X"FE",X"FC",X"FF",X"FC",X"FF",X"FE",X"FE",X"FF",X"FE",X"FF",X"FC",X"FC",X"FF",
		X"FD",X"FC",X"FE",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FD",X"FD",X"FC",X"FC",X"FD",X"FD",X"FF",
		X"FC",X"FE",X"FD",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FC",X"FE",X"FD",X"FE",X"FC",X"FE",X"FD",
		X"FE",X"FC",X"FC",X"FF",X"FE",X"FC",X"FD",X"FC",X"FD",X"FC",X"FC",X"FF",X"FC",X"FE",X"FC",X"FC",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FD",X"FC",X"FF",X"FD",X"FD",X"FF",X"FC",X"FF",X"FD",X"FC",X"FF",
		X"FD",X"FC",X"FD",X"FC",X"FD",X"FD",X"FD",X"FE",X"FD",X"FF",X"FD",X"FE",X"FE",X"FF",X"FE",X"FE",
		X"FF",X"FC",X"FD",X"FC",X"FF",X"FD",X"FC",X"FF",X"FF",X"FD",X"FE",X"FC",X"FD",X"FC",X"FD",X"FC",
		X"FD",X"FD",X"FD",X"FE",X"FC",X"FE",X"FC",X"FF",X"FF",X"FE",X"FE",X"FF",X"FD",X"FC",X"FE",X"FC",
		X"FF",X"FC",X"FF",X"FD",X"FF",X"FD",X"FD",X"FE",X"FE",X"FC",X"FD",X"FD",X"FC",X"FC",X"FC",X"FF",
		X"FD",X"FF",X"FC",X"FD",X"FF",X"FF",X"FE",X"FE",X"FF",X"FC",X"FC",X"FF",X"FC",X"FD",X"FC",X"FF",
		X"FF",X"FC",X"FD",X"FF",X"FD",X"FC",X"FC",X"FD",X"FC",X"FC",X"FD",X"FE",X"FD",X"FF",X"FC",X"FC",
		X"FE",X"FF",X"FE",X"FF",X"FF",X"FD",X"FF",X"FC",X"FD",X"FD",X"FE",X"FD",X"FD",X"FC",X"FD",X"FE",
		X"FF",X"FD",X"FC",X"FC",X"FD",X"FD",X"FD",X"FE",X"FC",X"FF",X"FC",X"FC",X"FF",X"FE",X"FF",X"FE",
		X"FF",X"FD",X"FC",X"FF",X"FD",X"FD",X"FE",X"FC",X"FC",X"FD",X"FD",X"FE",X"FD",X"FD",X"FD",X"FC",
		X"FC",X"FD",X"FD",X"FE",X"FC",X"FE",X"FC",X"FD",X"FF",X"FE",X"FE",X"FE",X"FF",X"FC",X"FD",X"FD",
		X"FF",X"FD",X"FD",X"FE",X"FE",X"FC",X"FF",X"FC",X"FD",X"FD",X"FC",X"FD",X"FD",X"FC",X"FC",X"FF",
		X"FD",X"FE",X"FC",X"FC",X"FF",X"FE",X"FE",X"FF",X"FC",X"FD",X"FC",X"FF",X"FF",X"FC",X"FF",X"FD",
		X"FD",X"FC",X"FC",X"FF",X"FF",X"FD",X"FD",X"FC",X"FC",X"FD",X"FD",X"FE",X"FC",X"FE",X"FD",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",
		X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FF",X"FD",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FD",X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FF",X"FD",X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FF",X"FD",X"FF",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FF",X"FD",
		X"FF",X"FF",X"FD",X"FD",X"FD",X"FF",X"FF",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FD",X"FF",X"FF",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FD",X"FF",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",
		X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FD",X"FD",X"FF",X"FD",X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FD",
		X"FF",X"FD",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AE");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
